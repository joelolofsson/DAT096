------------------------------------------------------------------------------
--  This file is a part of the GRLIB VHDL IP LIBRARY
--  Copyright (C) 2011, Aeroflex Gaisler AB - all rights reserved.
--
-- ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN 
-- ACCORDANCE WITH THE GAISLER LICENSE AGREEMENT AND MUST BE APPROVED 
-- IN ADVANCE IN WRITING. 
------------------------------------------------------------------------------
--
-- Written by Synplicity
-- Product Version "E-2010.09"
-- Program "Synplify Pro", Mapper "maprc, Build 140R"
-- Mon Jan 31 15:45:53 2011
--

--
-- Written by Synplify Pro version Build 140R
-- Mon Jan 31 15:45:53 2011
--

--
library ieee, stratixii;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
--library synplify;
--use synplify.components.all;
use stratixii.stratixii_components.all;

entity grlfpw_0_stratixii is
port(
  rst :  in std_logic;
  clk :  in std_logic;
  holdn :  in std_logic;
  cpi_flush :  in std_logic;
  cpi_exack :  in std_logic;
  cpi_a_rs1 : in std_logic_vector(4 downto 0);
  cpi_d_pc : in std_logic_vector(31 downto 0);
  cpi_d_inst : in std_logic_vector(31 downto 0);
  cpi_d_cnt : in std_logic_vector(1 downto 0);
  cpi_d_trap :  in std_logic;
  cpi_d_annul :  in std_logic;
  cpi_d_pv :  in std_logic;
  cpi_a_pc : in std_logic_vector(31 downto 0);
  cpi_a_inst : in std_logic_vector(31 downto 0);
  cpi_a_cnt : in std_logic_vector(1 downto 0);
  cpi_a_trap :  in std_logic;
  cpi_a_annul :  in std_logic;
  cpi_a_pv :  in std_logic;
  cpi_e_pc : in std_logic_vector(31 downto 0);
  cpi_e_inst : in std_logic_vector(31 downto 0);
  cpi_e_cnt : in std_logic_vector(1 downto 0);
  cpi_e_trap :  in std_logic;
  cpi_e_annul :  in std_logic;
  cpi_e_pv :  in std_logic;
  cpi_m_pc : in std_logic_vector(31 downto 0);
  cpi_m_inst : in std_logic_vector(31 downto 0);
  cpi_m_cnt : in std_logic_vector(1 downto 0);
  cpi_m_trap :  in std_logic;
  cpi_m_annul :  in std_logic;
  cpi_m_pv :  in std_logic;
  cpi_x_pc : in std_logic_vector(31 downto 0);
  cpi_x_inst : in std_logic_vector(31 downto 0);
  cpi_x_cnt : in std_logic_vector(1 downto 0);
  cpi_x_trap :  in std_logic;
  cpi_x_annul :  in std_logic;
  cpi_x_pv :  in std_logic;
  cpi_lddata : in std_logic_vector(31 downto 0);
  cpi_dbg_enable :  in std_logic;
  cpi_dbg_write :  in std_logic;
  cpi_dbg_fsr :  in std_logic;
  cpi_dbg_addr : in std_logic_vector(4 downto 0);
  cpi_dbg_data : in std_logic_vector(31 downto 0);
  cpo_data : out std_logic_vector(31 downto 0);
  cpo_exc :  out std_logic;
  cpo_cc : out std_logic_vector(1 downto 0);
  cpo_ccv :  out std_logic;
  cpo_ldlock :  out std_logic;
  cpo_holdn :  out std_logic;
  cpo_dbg_data : out std_logic_vector(31 downto 0);
  rfi1_rd1addr : out std_logic_vector(3 downto 0);
  rfi1_rd2addr : out std_logic_vector(3 downto 0);
  rfi1_wraddr : out std_logic_vector(3 downto 0);
  rfi1_wrdata : out std_logic_vector(31 downto 0);
  rfi1_ren1 :  out std_logic;
  rfi1_ren2 :  out std_logic;
  rfi1_wren :  out std_logic;
  rfi2_rd1addr : out std_logic_vector(3 downto 0);
  rfi2_rd2addr : out std_logic_vector(3 downto 0);
  rfi2_wraddr : out std_logic_vector(3 downto 0);
  rfi2_wrdata : out std_logic_vector(31 downto 0);
  rfi2_ren1 :  out std_logic;
  rfi2_ren2 :  out std_logic;
  rfi2_wren :  out std_logic;
  rfo1_data1 : in std_logic_vector(31 downto 0);
  rfo1_data2 : in std_logic_vector(31 downto 0);
  rfo2_data1 : in std_logic_vector(31 downto 0);
  rfo2_data2 : in std_logic_vector(31 downto 0));
end grlfpw_0_stratixii;

architecture beh of grlfpw_0_stratixii is
  signal devclrn : std_logic := '1';
  signal devpor : std_logic := '1';
  signal devoe : std_logic := '0';
  signal \GRLFPC2_0.FPI.OP2\ : std_logic_vector(63 downto 32);
  signal \GRLFPC2_0.R.FSR.RD\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.FPO.FRAC\ : std_logic_vector(54 downto 3);
  signal \GRLFPC2_0.FPO.EXP\ : std_logic_vector(10 downto 0);
  signal \GRLFPC2_0.R.STATE\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.R.I.INST\ : std_logic_vector(31 downto 0);
  signal \GRLFPC2_0.R.FSR.TEM\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.R.I.EXC\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.R.FSR.AEXC\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.R.A.RS1\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.R.A.RS2\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.R.FSR.CEXC\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.R.FSR.FTT\ : std_logic_vector(2 downto 0);
  signal \GRLFPC2_0.R.I.RES\ : std_logic_vector(63 downto 0);
  signal \GRLFPC2_0.COMB.V.I.RES_1\ : std_logic_vector(63 to 63);
  signal \GRLFPC2_0.R.A.RF1REN\ : std_logic_vector(2 downto 1);
  signal \GRLFPC2_0.R.A.RF2REN\ : std_logic_vector(2 downto 1);
  signal \GRLFPC2_0.FPCI_O_3\ : std_logic_vector(74 downto 0);
  signal \GRLFPC2_0.R.STATE_O_3\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.FPCI_O_0\ : std_logic_vector(70 downto 59);
  signal \GRLFPC2_0.FPCI_O\ : std_logic_vector(314 downto 0);
  signal \GRLFPC2_0.R.STATE_O\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.R.I.CC\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.R.I.PC_O\ : std_logic_vector(31 downto 2);
  signal \GRLFPC2_0.R.I.EXC_MB\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.COMB.RS1_1\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.COMB.RS2_1\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\ : std_logic_vector(85 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\ : std_logic_vector(16 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\ : std_logic_vector(377 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\ : std_logic_vector(57 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\ : std_logic_vector(12 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_57\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_56\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_55\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_54\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_53\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_52\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_51\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_50\ : std_logic_vector(7 to 7);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_49\ : std_logic_vector(8 to 8);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_48\ : std_logic_vector(9 to 9);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_47\ : std_logic_vector(10 to 10);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_46\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_45\ : std_logic_vector(12 to 12);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_44\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_43\ : std_logic_vector(14 to 14);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_42\ : std_logic_vector(15 to 15);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_41\ : std_logic_vector(16 to 16);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_40\ : std_logic_vector(17 to 17);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_39\ : std_logic_vector(18 to 18);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_38\ : std_logic_vector(19 to 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_37\ : std_logic_vector(20 to 20);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_36\ : std_logic_vector(21 to 21);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_35\ : std_logic_vector(22 to 22);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_34\ : std_logic_vector(23 to 23);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_33\ : std_logic_vector(24 to 24);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_32\ : std_logic_vector(25 to 25);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_31\ : std_logic_vector(26 to 26);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_30\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_29\ : std_logic_vector(28 to 28);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_28\ : std_logic_vector(29 to 29);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_27\ : std_logic_vector(30 to 30);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_26\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_25\ : std_logic_vector(32 to 32);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_24\ : std_logic_vector(33 to 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_23\ : std_logic_vector(34 to 34);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_22\ : std_logic_vector(35 to 35);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_21\ : std_logic_vector(36 to 36);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_20\ : std_logic_vector(37 to 37);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_19\ : std_logic_vector(38 to 38);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_18\ : std_logic_vector(39 to 39);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_17\ : std_logic_vector(40 to 40);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_16\ : std_logic_vector(41 to 41);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_15\ : std_logic_vector(42 to 42);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_14\ : std_logic_vector(43 to 43);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_13\ : std_logic_vector(44 to 44);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_12\ : std_logic_vector(45 to 45);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_11\ : std_logic_vector(46 to 46);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_10\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_9\ : std_logic_vector(48 to 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_8\ : std_logic_vector(49 to 49);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_7\ : std_logic_vector(50 to 50);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_6\ : std_logic_vector(51 to 51);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_5\ : std_logic_vector(52 to 52);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_113\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SBLSBS_1\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_112\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_111\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_110\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_109\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_108\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_107\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_106\ : std_logic_vector(7 to 7);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_105\ : std_logic_vector(8 to 8);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_104\ : std_logic_vector(9 to 9);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_103\ : std_logic_vector(10 to 10);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_102\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_101\ : std_logic_vector(12 to 12);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_100\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_99\ : std_logic_vector(14 to 14);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_98\ : std_logic_vector(15 to 15);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_97\ : std_logic_vector(16 to 16);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_96\ : std_logic_vector(17 to 17);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_95\ : std_logic_vector(18 to 18);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_94\ : std_logic_vector(19 to 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_93\ : std_logic_vector(20 to 20);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_92\ : std_logic_vector(21 to 21);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_91\ : std_logic_vector(22 to 22);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_90\ : std_logic_vector(23 to 23);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_89\ : std_logic_vector(24 to 24);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_88\ : std_logic_vector(25 to 25);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_87\ : std_logic_vector(26 to 26);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_86\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_85\ : std_logic_vector(28 to 28);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_84\ : std_logic_vector(29 to 29);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_83\ : std_logic_vector(30 to 30);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_82\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_81\ : std_logic_vector(32 to 32);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_80\ : std_logic_vector(33 to 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_79\ : std_logic_vector(34 to 34);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_78\ : std_logic_vector(35 to 35);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_77\ : std_logic_vector(36 to 36);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_76\ : std_logic_vector(37 to 37);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_75\ : std_logic_vector(38 to 38);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_74\ : std_logic_vector(39 to 39);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_73\ : std_logic_vector(40 to 40);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_72\ : std_logic_vector(41 to 41);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_71\ : std_logic_vector(42 to 42);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_70\ : std_logic_vector(43 to 43);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_69\ : std_logic_vector(44 to 44);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_68\ : std_logic_vector(45 to 45);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_67\ : std_logic_vector(46 to 46);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_66\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_65\ : std_logic_vector(48 to 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_64\ : std_logic_vector(49 to 49);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_63\ : std_logic_vector(50 to 50);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_62\ : std_logic_vector(51 to 51);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\ : std_logic_vector(57 downto 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SCLSBS_2\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SCLSBS_1\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_168\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_167\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_166\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_165\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_164\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_163\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_162\ : std_logic_vector(7 to 7);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_161\ : std_logic_vector(8 to 8);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_160\ : std_logic_vector(9 to 9);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_159\ : std_logic_vector(10 to 10);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_158\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_157\ : std_logic_vector(12 to 12);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_156\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_155\ : std_logic_vector(14 to 14);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_154\ : std_logic_vector(15 to 15);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_153\ : std_logic_vector(16 to 16);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_152\ : std_logic_vector(17 to 17);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_151\ : std_logic_vector(18 to 18);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_150\ : std_logic_vector(19 to 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_149\ : std_logic_vector(20 to 20);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_148\ : std_logic_vector(21 to 21);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_147\ : std_logic_vector(22 to 22);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_146\ : std_logic_vector(23 to 23);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_145\ : std_logic_vector(24 to 24);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_144\ : std_logic_vector(25 to 25);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_143\ : std_logic_vector(26 to 26);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_142\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_141\ : std_logic_vector(28 to 28);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_140\ : std_logic_vector(29 to 29);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_139\ : std_logic_vector(30 to 30);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_138\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_137\ : std_logic_vector(32 to 32);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_136\ : std_logic_vector(33 to 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_135\ : std_logic_vector(34 to 34);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_134\ : std_logic_vector(35 to 35);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_133\ : std_logic_vector(36 to 36);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_132\ : std_logic_vector(37 to 37);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_131\ : std_logic_vector(38 to 38);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_130\ : std_logic_vector(39 to 39);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_129\ : std_logic_vector(40 to 40);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_128\ : std_logic_vector(41 to 41);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_127\ : std_logic_vector(42 to 42);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_126\ : std_logic_vector(43 to 43);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_125\ : std_logic_vector(44 to 44);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_124\ : std_logic_vector(45 to 45);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_123\ : std_logic_vector(46 to 46);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_122\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_121\ : std_logic_vector(48 to 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_120\ : std_logic_vector(49 to 49);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_119\ : std_logic_vector(50 to 50);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\ : std_logic_vector(55 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\ : std_logic_vector(112 downto 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\ : std_logic_vector(9 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\ : std_logic_vector(2 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\ : std_logic_vector(12 downto 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_DIVMULTV\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\ : std_logic_vector(375 downto 58);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_14\ : std_logic_vector(172 downto 142);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\ : std_logic_vector(112 downto 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SCTRL_NEW\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW_6\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19\ : std_logic_vector(45 downto 9);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\ : std_logic_vector(112 downto 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M\ : std_logic_vector(6 downto 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT\ : std_logic_vector(4 downto 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M\ : std_logic_vector(79 to 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M\ : std_logic_vector(84 to 84);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_5\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_1\ : std_logic_vector(30 to 30);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_58\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.FPI.OP1\ : std_logic_vector(63 downto 32);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\ : std_logic_vector(8 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\ : std_logic_vector(4 downto 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SALSBS_1\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SALSBS_2\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M2\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12\ : std_logic_vector(2 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M13\ : std_logic_vector(2 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M8\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\ : std_logic_vector(54 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\ : std_logic_vector(57 downto 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\ : std_logic_vector(113 downto 58);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\ : std_logic_vector(8 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\ : std_logic_vector(9 downto 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.R.I.PC\ : std_logic_vector(30 downto 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_41\ : std_logic_vector(255 downto 251);
  signal \GRLFPC2_0.COMB.V.A.RF2REN_1_1\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.COMB.WRDATA_4\ : std_logic_vector(62 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\ : std_logic_vector(115 downto 114);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\ : std_logic_vector(115 downto 114);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\ : std_logic_vector(55 downto 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\ : std_logic_vector(18 downto 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.U_RDN_1\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\ : std_logic_vector(54 downto 15);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\ : std_logic_vector(56 downto 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\ : std_logic_vector(6 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\ : std_logic_vector(56 downto 46);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\ : std_logic_vector(5 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8_0\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SBLSBS_2\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_8_0\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_4\ : std_logic_vector(47 downto 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_13_C\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_9_TZ\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_22_1\ : std_logic_vector(52 to 52);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_4_0\ : std_logic_vector(34 to 34);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_6_1\ : std_logic_vector(25 to 25);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_6_1\ : std_logic_vector(58 to 58);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_11_1\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A9_3_0\ : std_logic_vector(28 to 28);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_9_0\ : std_logic_vector(62 downto 50);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_I_I_0\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_3_I\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\ : std_logic_vector(57 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\ : std_logic_vector(55 downto 46);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\ : std_logic_vector(49 downto 9);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\ : std_logic_vector(45 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_I_0_A2_4\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_4\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_6\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_7_1\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_1_1\ : std_logic_vector(58 to 58);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_25_1\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A24_8_1\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_A26_6_1\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_15_0\ : std_logic_vector(58 to 58);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_A26_23_0\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_44_0\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_3_0\ : std_logic_vector(18 to 18);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_2_0\ : std_logic_vector(58 to 58);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_31_1\ : std_logic_vector(48 to 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A24_10_1\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_13_0\ : std_logic_vector(59 to 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A24_1_0\ : std_logic_vector(55 downto 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_19_1\ : std_logic_vector(53 to 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_2_0\ : std_logic_vector(17 to 17);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A24_17_0\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O27_1_0\ : std_logic_vector(58 to 58);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_9_1\ : std_logic_vector(50 to 50);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_39_0\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_9_0\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_38_0\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2_1\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_5_2\ : std_logic_vector(52 to 52);
  signal \GRLFPC2_0.R.FSR.FTT_M_2\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_7_0\ : std_logic_vector(52 to 52);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A28_24_0\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_24_3\ : std_logic_vector(32 to 32);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_10_3\ : std_logic_vector(59 to 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A28_0_0\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A9_0_1\ : std_logic_vector(28 to 28);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_22_0\ : std_logic_vector(52 to 52);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_11_0\ : std_logic_vector(49 to 49);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_6_1\ : std_logic_vector(53 to 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_12_0\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A12_0_0\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_A26_7_0\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_3_0\ : std_logic_vector(25 to 25);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A21_0\ : std_logic_vector(59 to 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_0_0\ : std_logic_vector(17 to 17);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4_0\ : std_logic_vector(59 to 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A12_0\ : std_logic_vector(61 to 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_25_0\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_6_0\ : std_logic_vector(52 to 52);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3_0\ : std_logic_vector(41 to 41);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_22_0\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_20_0\ : std_logic_vector(7 to 7);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_9_0\ : std_logic_vector(19 to 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A3_0\ : std_logic_vector(26 to 26);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0_0\ : std_logic_vector(34 to 34);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_15_0\ : std_logic_vector(7 to 7);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A17_0\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_13_0\ : std_logic_vector(36 to 36);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_6_2\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_6_3\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_1_0\ : std_logic_vector(39 to 39);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O2_1\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O2_2\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_0\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_1\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_3\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_5\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_6\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_7\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_9_0\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_10\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_12\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_15_0\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_19\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_21\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_23\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_0\ : std_logic_vector(47 downto 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_2\ : std_logic_vector(47 downto 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_3\ : std_logic_vector(47 downto 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_5\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_8\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_9\ : std_logic_vector(47 downto 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_10\ : std_logic_vector(47 downto 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_12\ : std_logic_vector(47 downto 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_13\ : std_logic_vector(47 downto 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_14\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_20\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_1_2\ : std_logic_vector(22 to 22);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_6\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_15\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_17\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_22\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_23\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV_0\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0\ : std_logic_vector(9 to 9);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_IV_0\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_4_0\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_4_0\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8_I\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\ : std_logic_vector(15 downto 8);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\ : std_logic_vector(231 downto 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_5_2_RETO\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\ : std_logic_vector(84 downto 49);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO\ : std_logic_vector(1 to 1);
  signal CPI_D_INST_RETO : std_logic_vector(12 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO\ : std_logic_vector(2 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO\ : std_logic_vector(6 downto 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO\ : std_logic_vector(55 downto 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO\ : std_logic_vector(79 to 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO\ : std_logic_vector(84 to 84);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_4_0_RETO\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_2_RETO\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_5_1_RETO\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_I_I_0_RETO\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.U_RDN_1_RETO\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_RETO\ : std_logic_vector(9 downto 8);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\ : std_logic_vector(99 downto 72);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\ : std_logic_vector(106 downto 68);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1_RETO\ : std_logic_vector(115 downto 72);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0_RETO\ : std_logic_vector(115 downto 72);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\ : std_logic_vector(106 downto 68);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\ : std_logic_vector(4 downto 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_3_I_RETO\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\ : std_logic_vector(113 downto 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_RETO\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0_RETO\ : std_logic_vector(9 to 9);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_RETO\ : std_logic_vector(12 to 12);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_13_C_RETO\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\ : std_logic_vector(98 downto 1);
  signal \GRLFPC2_0.FPO.FRAC_RETO\ : std_logic_vector(54 downto 15);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_4_0_RETO\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\ : std_logic_vector(73 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\ : std_logic_vector(73 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI_0\ : std_logic_vector(10 to 10);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_229\ : std_logic_vector(78 to 78);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\ : std_logic_vector(84 downto 81);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\ : std_logic_vector(84 downto 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\ : std_logic_vector(81 downto 78);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\ : std_logic_vector(81 downto 78);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\ : std_logic_vector(84 downto 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\ : std_logic_vector(84 downto 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\ : std_logic_vector(81 downto 78);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\ : std_logic_vector(8 downto 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\ : std_logic_vector(241 downto 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\ : std_logic_vector(8 downto 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\ : std_logic_vector(241 downto 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\ : std_logic_vector(3 downto 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_0\ : std_logic_vector(15 to 15);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\ : std_logic_vector(3 downto 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\ : std_logic_vector(43 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_1\ : std_logic_vector(15 to 15);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\ : std_logic_vector(43 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_2\ : std_logic_vector(15 to 15);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\ : std_logic_vector(42 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_3\ : std_logic_vector(15 to 15);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\ : std_logic_vector(3 downto 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_0\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\ : std_logic_vector(3 downto 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_1\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\ : std_logic_vector(57 downto 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2_0\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2_1\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\ : std_logic_vector(42 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_4\ : std_logic_vector(15 to 15);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_6\ : std_logic_vector(42 to 42);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_5\ : std_logic_vector(15 to 15);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_0\ : std_logic_vector(8 downto 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_3\ : std_logic_vector(55 downto 21);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_1\ : std_logic_vector(6 downto 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_4\ : std_logic_vector(53 downto 21);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19_0\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19_1\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_6\ : std_logic_vector(15 to 15);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_7\ : std_logic_vector(42 to 42);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\ : std_logic_vector(81 downto 78);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_0\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\ : std_logic_vector(81 to 81);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_1\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\ : std_logic_vector(81 to 81);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_2\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\ : std_logic_vector(81 to 81);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_3\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\ : std_logic_vector(81 to 81);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_4\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_5\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\ : std_logic_vector(84 downto 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_6\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\ : std_logic_vector(84 downto 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_7\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\ : std_logic_vector(84 downto 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_8\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\ : std_logic_vector(84 downto 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_9\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_0\ : std_logic_vector(1 to 1);
  signal CPI_D_INST_RETO_0 : std_logic_vector(12 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_1\ : std_logic_vector(1 to 1);
  signal CPI_D_INST_RETO_1 : std_logic_vector(12 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_2\ : std_logic_vector(1 to 1);
  signal CPI_D_INST_RETO_2 : std_logic_vector(12 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_3\ : std_logic_vector(1 to 1);
  signal CPI_D_INST_RETO_3 : std_logic_vector(12 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_4\ : std_logic_vector(1 to 1);
  signal CPI_D_INST_RETO_4 : std_logic_vector(12 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_5\ : std_logic_vector(1 to 1);
  signal CPI_D_INST_RETO_5 : std_logic_vector(12 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_6\ : std_logic_vector(1 to 1);
  signal CPI_D_INST_RETO_6 : std_logic_vector(12 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\ : std_logic_vector(84 downto 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_7\ : std_logic_vector(1 to 1);
  signal CPI_D_INST_RETO_7 : std_logic_vector(12 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\ : std_logic_vector(83 downto 82);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\ : std_logic_vector(82 downto 49);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\ : std_logic_vector(83 downto 82);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\ : std_logic_vector(82 downto 65);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\ : std_logic_vector(83 downto 82);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_2\ : std_logic_vector(82 to 82);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\ : std_logic_vector(83 downto 82);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_3\ : std_logic_vector(82 to 82);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\ : std_logic_vector(83 downto 82);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_4\ : std_logic_vector(82 to 82);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\ : std_logic_vector(83 downto 82);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_5\ : std_logic_vector(82 to 82);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\ : std_logic_vector(83 downto 82);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_6\ : std_logic_vector(82 to 82);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\ : std_logic_vector(82 to 82);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_7\ : std_logic_vector(82 to 82);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\ : std_logic_vector(82 to 82);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_8\ : std_logic_vector(82 to 82);
  signal CPI_D_INST_RETO_8 : std_logic_vector(12 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\ : std_logic_vector(83 to 83);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_0\ : std_logic_vector(2 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_0\ : std_logic_vector(6 downto 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\ : std_logic_vector(83 to 83);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_1\ : std_logic_vector(2 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_1\ : std_logic_vector(6 downto 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\ : std_logic_vector(83 to 83);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_2\ : std_logic_vector(2 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_2\ : std_logic_vector(6 downto 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_3\ : std_logic_vector(2 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_3\ : std_logic_vector(6 downto 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_4\ : std_logic_vector(2 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_4\ : std_logic_vector(6 downto 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_5\ : std_logic_vector(2 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_5\ : std_logic_vector(6 downto 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_6\ : std_logic_vector(2 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_6\ : std_logic_vector(6 downto 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_7\ : std_logic_vector(2 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_7\ : std_logic_vector(6 downto 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_8\ : std_logic_vector(2 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_8\ : std_logic_vector(6 downto 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_9\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_9\ : std_logic_vector(2 to 2);
  signal CPI_D_INST_RETO_9 : std_logic_vector(7 to 7);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\ : std_logic_vector(85 to 85);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\ : std_logic_vector(85 to 85);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\ : std_logic_vector(85 to 85);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\ : std_logic_vector(85 to 85);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\ : std_logic_vector(85 to 85);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\ : std_logic_vector(85 to 85);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\ : std_logic_vector(85 to 85);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\ : std_logic_vector(85 to 85);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\ : std_logic_vector(85 to 85);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_0\ : std_logic_vector(55 downto 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO_0\ : std_logic_vector(79 to 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\ : std_logic_vector(80 downto 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_1\ : std_logic_vector(55 downto 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO_1\ : std_logic_vector(79 to 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\ : std_logic_vector(80 to 80);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_2\ : std_logic_vector(55 downto 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO_2\ : std_logic_vector(79 to 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\ : std_logic_vector(80 to 80);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_3\ : std_logic_vector(55 downto 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO_3\ : std_logic_vector(79 to 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\ : std_logic_vector(80 to 80);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_4\ : std_logic_vector(55 downto 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO_4\ : std_logic_vector(79 to 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\ : std_logic_vector(80 to 80);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_5\ : std_logic_vector(55 downto 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO_5\ : std_logic_vector(79 to 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\ : std_logic_vector(80 to 80);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_6\ : std_logic_vector(55 downto 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO_6\ : std_logic_vector(79 to 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\ : std_logic_vector(80 to 80);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_7\ : std_logic_vector(55 downto 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO_7\ : std_logic_vector(79 to 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\ : std_logic_vector(80 to 80);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_8\ : std_logic_vector(55 downto 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO_8\ : std_logic_vector(79 to 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\ : std_logic_vector(78 to 78);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO_0\ : std_logic_vector(84 to 84);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\ : std_logic_vector(78 to 78);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO_1\ : std_logic_vector(84 to 84);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\ : std_logic_vector(78 to 78);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO_2\ : std_logic_vector(84 to 84);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\ : std_logic_vector(78 to 78);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO_3\ : std_logic_vector(84 to 84);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\ : std_logic_vector(78 to 78);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO_4\ : std_logic_vector(84 to 84);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO_5\ : std_logic_vector(84 to 84);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO_6\ : std_logic_vector(84 to 84);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO_7\ : std_logic_vector(84 to 84);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO_8\ : std_logic_vector(84 to 84);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251_0\ : std_logic_vector(80 to 80);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238_0\ : std_logic_vector(81 to 81);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_5\ : std_logic_vector(53 downto 21);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_6\ : std_logic_vector(53 downto 21);
  signal CPO_DATAZ : std_logic_vector(31 downto 0);
  signal CPO_CCZ : std_logic_vector(1 downto 0);
  signal CPO_DBG_DATAZ : std_logic_vector(31 downto 0);
  signal RFI1_WRDATAZ : std_logic_vector(31 downto 0);
  signal RFI2_RD1ADDRZ : std_logic_vector(3 downto 0);
  signal RFI2_RD2ADDRZ : std_logic_vector(3 downto 0);
  signal RFI2_WRADDRZ : std_logic_vector(3 downto 0);
  signal RFI2_WRDATAZ : std_logic_vector(31 downto 0);
  signal CLK_INTERNAL : std_logic ;
  signal HOLDN_INTERNAL : std_logic ;
  signal CPI_FLUSH_INTERNAL : std_logic ;
  signal CPI_EXACK_INTERNAL : std_logic ;
  signal CPI_A_RS1_INTERNAL : std_logic ;
  signal CPI_A_RS1_INTERNAL_0 : std_logic ;
  signal CPI_A_RS1_INTERNAL_1 : std_logic ;
  signal CPI_A_RS1_INTERNAL_2 : std_logic ;
  signal CPI_A_RS1_INTERNAL_3 : std_logic ;
  signal CPI_D_PC_INTERNAL : std_logic ;
  signal CPI_D_PC_INTERNAL_0 : std_logic ;
  signal CPI_D_PC_INTERNAL_1 : std_logic ;
  signal CPI_D_PC_INTERNAL_2 : std_logic ;
  signal CPI_D_PC_INTERNAL_3 : std_logic ;
  signal CPI_D_PC_INTERNAL_4 : std_logic ;
  signal CPI_D_PC_INTERNAL_5 : std_logic ;
  signal CPI_D_PC_INTERNAL_6 : std_logic ;
  signal CPI_D_PC_INTERNAL_7 : std_logic ;
  signal CPI_D_PC_INTERNAL_8 : std_logic ;
  signal CPI_D_PC_INTERNAL_9 : std_logic ;
  signal CPI_D_PC_INTERNAL_10 : std_logic ;
  signal CPI_D_PC_INTERNAL_11 : std_logic ;
  signal CPI_D_PC_INTERNAL_12 : std_logic ;
  signal CPI_D_PC_INTERNAL_13 : std_logic ;
  signal CPI_D_PC_INTERNAL_14 : std_logic ;
  signal CPI_D_PC_INTERNAL_15 : std_logic ;
  signal CPI_D_PC_INTERNAL_16 : std_logic ;
  signal CPI_D_PC_INTERNAL_17 : std_logic ;
  signal CPI_D_PC_INTERNAL_18 : std_logic ;
  signal CPI_D_PC_INTERNAL_19 : std_logic ;
  signal CPI_D_PC_INTERNAL_20 : std_logic ;
  signal CPI_D_PC_INTERNAL_21 : std_logic ;
  signal CPI_D_PC_INTERNAL_22 : std_logic ;
  signal CPI_D_PC_INTERNAL_23 : std_logic ;
  signal CPI_D_PC_INTERNAL_24 : std_logic ;
  signal CPI_D_PC_INTERNAL_25 : std_logic ;
  signal CPI_D_PC_INTERNAL_26 : std_logic ;
  signal CPI_D_PC_INTERNAL_27 : std_logic ;
  signal CPI_D_PC_INTERNAL_28 : std_logic ;
  signal CPI_D_PC_INTERNAL_29 : std_logic ;
  signal CPI_D_PC_INTERNAL_30 : std_logic ;
  signal CPI_D_INST_INTERNAL : std_logic ;
  signal CPI_D_INST_INTERNAL_0 : std_logic ;
  signal CPI_D_INST_INTERNAL_1 : std_logic ;
  signal CPI_D_INST_INTERNAL_2 : std_logic ;
  signal CPI_D_INST_INTERNAL_3 : std_logic ;
  signal CPI_D_INST_INTERNAL_4 : std_logic ;
  signal CPI_D_INST_INTERNAL_5 : std_logic ;
  signal CPI_D_INST_INTERNAL_7 : std_logic ;
  signal CPI_D_INST_INTERNAL_8 : std_logic ;
  signal CPI_D_INST_INTERNAL_9 : std_logic ;
  signal CPI_D_INST_INTERNAL_10 : std_logic ;
  signal CPI_D_INST_INTERNAL_11 : std_logic ;
  signal CPI_D_INST_INTERNAL_12 : std_logic ;
  signal CPI_D_INST_INTERNAL_13 : std_logic ;
  signal CPI_D_INST_INTERNAL_14 : std_logic ;
  signal CPI_D_INST_INTERNAL_15 : std_logic ;
  signal CPI_D_INST_INTERNAL_16 : std_logic ;
  signal CPI_D_INST_INTERNAL_17 : std_logic ;
  signal CPI_D_INST_INTERNAL_18 : std_logic ;
  signal CPI_D_INST_INTERNAL_19 : std_logic ;
  signal CPI_D_INST_INTERNAL_20 : std_logic ;
  signal CPI_D_INST_INTERNAL_21 : std_logic ;
  signal CPI_D_INST_INTERNAL_22 : std_logic ;
  signal CPI_D_INST_INTERNAL_23 : std_logic ;
  signal CPI_D_INST_INTERNAL_24 : std_logic ;
  signal CPI_D_INST_INTERNAL_25 : std_logic ;
  signal CPI_D_INST_INTERNAL_26 : std_logic ;
  signal CPI_D_INST_INTERNAL_27 : std_logic ;
  signal CPI_D_INST_INTERNAL_28 : std_logic ;
  signal CPI_D_INST_INTERNAL_29 : std_logic ;
  signal CPI_D_INST_INTERNAL_30 : std_logic ;
  signal CPI_D_CNT_INTERNAL : std_logic ;
  signal CPI_D_CNT_INTERNAL_0 : std_logic ;
  signal CPI_D_TRAP_INTERNAL : std_logic ;
  signal CPI_D_ANNUL_INTERNAL : std_logic ;
  signal CPI_D_PV_INTERNAL : std_logic ;
  signal CPI_A_PC_INTERNAL : std_logic ;
  signal CPI_A_PC_INTERNAL_0 : std_logic ;
  signal CPI_A_PC_INTERNAL_1 : std_logic ;
  signal CPI_A_PC_INTERNAL_2 : std_logic ;
  signal CPI_A_PC_INTERNAL_3 : std_logic ;
  signal CPI_A_PC_INTERNAL_4 : std_logic ;
  signal CPI_A_PC_INTERNAL_5 : std_logic ;
  signal CPI_A_PC_INTERNAL_6 : std_logic ;
  signal CPI_A_PC_INTERNAL_7 : std_logic ;
  signal CPI_A_PC_INTERNAL_8 : std_logic ;
  signal CPI_A_PC_INTERNAL_9 : std_logic ;
  signal CPI_A_PC_INTERNAL_10 : std_logic ;
  signal CPI_A_PC_INTERNAL_11 : std_logic ;
  signal CPI_A_PC_INTERNAL_12 : std_logic ;
  signal CPI_A_PC_INTERNAL_13 : std_logic ;
  signal CPI_A_PC_INTERNAL_14 : std_logic ;
  signal CPI_A_PC_INTERNAL_15 : std_logic ;
  signal CPI_A_PC_INTERNAL_16 : std_logic ;
  signal CPI_A_PC_INTERNAL_17 : std_logic ;
  signal CPI_A_PC_INTERNAL_18 : std_logic ;
  signal CPI_A_PC_INTERNAL_19 : std_logic ;
  signal CPI_A_PC_INTERNAL_20 : std_logic ;
  signal CPI_A_PC_INTERNAL_21 : std_logic ;
  signal CPI_A_PC_INTERNAL_22 : std_logic ;
  signal CPI_A_PC_INTERNAL_23 : std_logic ;
  signal CPI_A_PC_INTERNAL_24 : std_logic ;
  signal CPI_A_PC_INTERNAL_25 : std_logic ;
  signal CPI_A_PC_INTERNAL_26 : std_logic ;
  signal CPI_A_PC_INTERNAL_27 : std_logic ;
  signal CPI_A_PC_INTERNAL_28 : std_logic ;
  signal CPI_A_PC_INTERNAL_29 : std_logic ;
  signal CPI_A_PC_INTERNAL_30 : std_logic ;
  signal CPI_A_INST_INTERNAL : std_logic ;
  signal CPI_A_INST_INTERNAL_0 : std_logic ;
  signal CPI_A_INST_INTERNAL_1 : std_logic ;
  signal CPI_A_INST_INTERNAL_2 : std_logic ;
  signal CPI_A_INST_INTERNAL_3 : std_logic ;
  signal CPI_A_INST_INTERNAL_4 : std_logic ;
  signal CPI_A_INST_INTERNAL_5 : std_logic ;
  signal CPI_A_INST_INTERNAL_6 : std_logic ;
  signal CPI_A_INST_INTERNAL_7 : std_logic ;
  signal CPI_A_INST_INTERNAL_8 : std_logic ;
  signal CPI_A_INST_INTERNAL_9 : std_logic ;
  signal CPI_A_INST_INTERNAL_10 : std_logic ;
  signal CPI_A_INST_INTERNAL_11 : std_logic ;
  signal CPI_A_INST_INTERNAL_12 : std_logic ;
  signal CPI_A_INST_INTERNAL_13 : std_logic ;
  signal CPI_A_INST_INTERNAL_14 : std_logic ;
  signal CPI_A_INST_INTERNAL_15 : std_logic ;
  signal CPI_A_INST_INTERNAL_16 : std_logic ;
  signal CPI_A_INST_INTERNAL_17 : std_logic ;
  signal CPI_A_INST_INTERNAL_18 : std_logic ;
  signal CPI_A_INST_INTERNAL_19 : std_logic ;
  signal CPI_A_INST_INTERNAL_20 : std_logic ;
  signal CPI_A_INST_INTERNAL_21 : std_logic ;
  signal CPI_A_INST_INTERNAL_22 : std_logic ;
  signal CPI_A_INST_INTERNAL_23 : std_logic ;
  signal CPI_A_INST_INTERNAL_24 : std_logic ;
  signal CPI_A_INST_INTERNAL_25 : std_logic ;
  signal CPI_A_INST_INTERNAL_26 : std_logic ;
  signal CPI_A_INST_INTERNAL_27 : std_logic ;
  signal CPI_A_INST_INTERNAL_28 : std_logic ;
  signal CPI_A_INST_INTERNAL_29 : std_logic ;
  signal CPI_A_INST_INTERNAL_30 : std_logic ;
  signal CPI_A_CNT_INTERNAL : std_logic ;
  signal CPI_A_CNT_INTERNAL_0 : std_logic ;
  signal CPI_A_TRAP_INTERNAL : std_logic ;
  signal CPI_A_ANNUL_INTERNAL : std_logic ;
  signal CPI_A_PV_INTERNAL : std_logic ;
  signal CPI_E_PC_INTERNAL : std_logic ;
  signal CPI_E_PC_INTERNAL_0 : std_logic ;
  signal CPI_E_PC_INTERNAL_1 : std_logic ;
  signal CPI_E_PC_INTERNAL_2 : std_logic ;
  signal CPI_E_PC_INTERNAL_3 : std_logic ;
  signal CPI_E_PC_INTERNAL_4 : std_logic ;
  signal CPI_E_PC_INTERNAL_5 : std_logic ;
  signal CPI_E_PC_INTERNAL_6 : std_logic ;
  signal CPI_E_PC_INTERNAL_7 : std_logic ;
  signal CPI_E_PC_INTERNAL_8 : std_logic ;
  signal CPI_E_PC_INTERNAL_9 : std_logic ;
  signal CPI_E_PC_INTERNAL_10 : std_logic ;
  signal CPI_E_PC_INTERNAL_11 : std_logic ;
  signal CPI_E_PC_INTERNAL_12 : std_logic ;
  signal CPI_E_PC_INTERNAL_13 : std_logic ;
  signal CPI_E_PC_INTERNAL_14 : std_logic ;
  signal CPI_E_PC_INTERNAL_15 : std_logic ;
  signal CPI_E_PC_INTERNAL_16 : std_logic ;
  signal CPI_E_PC_INTERNAL_17 : std_logic ;
  signal CPI_E_PC_INTERNAL_18 : std_logic ;
  signal CPI_E_PC_INTERNAL_19 : std_logic ;
  signal CPI_E_PC_INTERNAL_20 : std_logic ;
  signal CPI_E_PC_INTERNAL_21 : std_logic ;
  signal CPI_E_PC_INTERNAL_22 : std_logic ;
  signal CPI_E_PC_INTERNAL_23 : std_logic ;
  signal CPI_E_PC_INTERNAL_24 : std_logic ;
  signal CPI_E_PC_INTERNAL_25 : std_logic ;
  signal CPI_E_PC_INTERNAL_26 : std_logic ;
  signal CPI_E_PC_INTERNAL_27 : std_logic ;
  signal CPI_E_PC_INTERNAL_28 : std_logic ;
  signal CPI_E_PC_INTERNAL_29 : std_logic ;
  signal CPI_E_PC_INTERNAL_30 : std_logic ;
  signal CPI_E_INST_INTERNAL : std_logic ;
  signal CPI_E_INST_INTERNAL_0 : std_logic ;
  signal CPI_E_INST_INTERNAL_1 : std_logic ;
  signal CPI_E_INST_INTERNAL_2 : std_logic ;
  signal CPI_E_INST_INTERNAL_3 : std_logic ;
  signal CPI_E_INST_INTERNAL_4 : std_logic ;
  signal CPI_E_INST_INTERNAL_5 : std_logic ;
  signal CPI_E_INST_INTERNAL_6 : std_logic ;
  signal CPI_E_INST_INTERNAL_7 : std_logic ;
  signal CPI_E_INST_INTERNAL_8 : std_logic ;
  signal CPI_E_INST_INTERNAL_9 : std_logic ;
  signal CPI_E_INST_INTERNAL_10 : std_logic ;
  signal CPI_E_INST_INTERNAL_11 : std_logic ;
  signal CPI_E_INST_INTERNAL_12 : std_logic ;
  signal CPI_E_INST_INTERNAL_13 : std_logic ;
  signal CPI_E_INST_INTERNAL_14 : std_logic ;
  signal CPI_E_INST_INTERNAL_15 : std_logic ;
  signal CPI_E_INST_INTERNAL_16 : std_logic ;
  signal CPI_E_INST_INTERNAL_17 : std_logic ;
  signal CPI_E_INST_INTERNAL_18 : std_logic ;
  signal CPI_E_INST_INTERNAL_19 : std_logic ;
  signal CPI_E_INST_INTERNAL_20 : std_logic ;
  signal CPI_E_INST_INTERNAL_21 : std_logic ;
  signal CPI_E_INST_INTERNAL_22 : std_logic ;
  signal CPI_E_INST_INTERNAL_23 : std_logic ;
  signal CPI_E_INST_INTERNAL_24 : std_logic ;
  signal CPI_E_INST_INTERNAL_25 : std_logic ;
  signal CPI_E_INST_INTERNAL_26 : std_logic ;
  signal CPI_E_INST_INTERNAL_27 : std_logic ;
  signal CPI_E_INST_INTERNAL_28 : std_logic ;
  signal CPI_E_INST_INTERNAL_29 : std_logic ;
  signal CPI_E_INST_INTERNAL_30 : std_logic ;
  signal CPI_E_CNT_INTERNAL : std_logic ;
  signal CPI_E_CNT_INTERNAL_0 : std_logic ;
  signal CPI_E_TRAP_INTERNAL : std_logic ;
  signal CPI_E_ANNUL_INTERNAL : std_logic ;
  signal CPI_E_PV_INTERNAL : std_logic ;
  signal CPI_M_PC_INTERNAL : std_logic ;
  signal CPI_M_PC_INTERNAL_0 : std_logic ;
  signal CPI_M_PC_INTERNAL_1 : std_logic ;
  signal CPI_M_PC_INTERNAL_2 : std_logic ;
  signal CPI_M_PC_INTERNAL_3 : std_logic ;
  signal CPI_M_PC_INTERNAL_4 : std_logic ;
  signal CPI_M_PC_INTERNAL_5 : std_logic ;
  signal CPI_M_PC_INTERNAL_6 : std_logic ;
  signal CPI_M_PC_INTERNAL_7 : std_logic ;
  signal CPI_M_PC_INTERNAL_8 : std_logic ;
  signal CPI_M_PC_INTERNAL_9 : std_logic ;
  signal CPI_M_PC_INTERNAL_10 : std_logic ;
  signal CPI_M_PC_INTERNAL_11 : std_logic ;
  signal CPI_M_PC_INTERNAL_12 : std_logic ;
  signal CPI_M_PC_INTERNAL_13 : std_logic ;
  signal CPI_M_PC_INTERNAL_14 : std_logic ;
  signal CPI_M_PC_INTERNAL_15 : std_logic ;
  signal CPI_M_PC_INTERNAL_16 : std_logic ;
  signal CPI_M_PC_INTERNAL_17 : std_logic ;
  signal CPI_M_PC_INTERNAL_18 : std_logic ;
  signal CPI_M_PC_INTERNAL_19 : std_logic ;
  signal CPI_M_PC_INTERNAL_20 : std_logic ;
  signal CPI_M_PC_INTERNAL_21 : std_logic ;
  signal CPI_M_PC_INTERNAL_22 : std_logic ;
  signal CPI_M_PC_INTERNAL_23 : std_logic ;
  signal CPI_M_PC_INTERNAL_24 : std_logic ;
  signal CPI_M_PC_INTERNAL_25 : std_logic ;
  signal CPI_M_PC_INTERNAL_26 : std_logic ;
  signal CPI_M_PC_INTERNAL_27 : std_logic ;
  signal CPI_M_PC_INTERNAL_28 : std_logic ;
  signal CPI_M_PC_INTERNAL_29 : std_logic ;
  signal CPI_M_PC_INTERNAL_30 : std_logic ;
  signal CPI_M_INST_INTERNAL : std_logic ;
  signal CPI_M_INST_INTERNAL_0 : std_logic ;
  signal CPI_M_INST_INTERNAL_1 : std_logic ;
  signal CPI_M_INST_INTERNAL_2 : std_logic ;
  signal CPI_M_INST_INTERNAL_3 : std_logic ;
  signal CPI_M_INST_INTERNAL_4 : std_logic ;
  signal CPI_M_INST_INTERNAL_5 : std_logic ;
  signal CPI_M_INST_INTERNAL_6 : std_logic ;
  signal CPI_M_INST_INTERNAL_7 : std_logic ;
  signal CPI_M_INST_INTERNAL_8 : std_logic ;
  signal CPI_M_INST_INTERNAL_9 : std_logic ;
  signal CPI_M_INST_INTERNAL_10 : std_logic ;
  signal CPI_M_INST_INTERNAL_11 : std_logic ;
  signal CPI_M_INST_INTERNAL_12 : std_logic ;
  signal CPI_M_INST_INTERNAL_13 : std_logic ;
  signal CPI_M_INST_INTERNAL_14 : std_logic ;
  signal CPI_M_INST_INTERNAL_15 : std_logic ;
  signal CPI_M_INST_INTERNAL_16 : std_logic ;
  signal CPI_M_INST_INTERNAL_17 : std_logic ;
  signal CPI_M_INST_INTERNAL_18 : std_logic ;
  signal CPI_M_INST_INTERNAL_19 : std_logic ;
  signal CPI_M_INST_INTERNAL_20 : std_logic ;
  signal CPI_M_INST_INTERNAL_21 : std_logic ;
  signal CPI_M_INST_INTERNAL_22 : std_logic ;
  signal CPI_M_INST_INTERNAL_23 : std_logic ;
  signal CPI_M_INST_INTERNAL_24 : std_logic ;
  signal CPI_M_INST_INTERNAL_25 : std_logic ;
  signal CPI_M_INST_INTERNAL_26 : std_logic ;
  signal CPI_M_INST_INTERNAL_27 : std_logic ;
  signal CPI_M_INST_INTERNAL_28 : std_logic ;
  signal CPI_M_INST_INTERNAL_29 : std_logic ;
  signal CPI_M_INST_INTERNAL_30 : std_logic ;
  signal CPI_M_CNT_INTERNAL : std_logic ;
  signal CPI_M_CNT_INTERNAL_0 : std_logic ;
  signal CPI_M_TRAP_INTERNAL : std_logic ;
  signal CPI_M_ANNUL_INTERNAL : std_logic ;
  signal CPI_M_PV_INTERNAL : std_logic ;
  signal CPI_X_PC_INTERNAL : std_logic ;
  signal CPI_X_PC_INTERNAL_0 : std_logic ;
  signal CPI_X_PC_INTERNAL_1 : std_logic ;
  signal CPI_X_PC_INTERNAL_2 : std_logic ;
  signal CPI_X_PC_INTERNAL_3 : std_logic ;
  signal CPI_X_PC_INTERNAL_4 : std_logic ;
  signal CPI_X_PC_INTERNAL_5 : std_logic ;
  signal CPI_X_PC_INTERNAL_6 : std_logic ;
  signal CPI_X_PC_INTERNAL_7 : std_logic ;
  signal CPI_X_PC_INTERNAL_8 : std_logic ;
  signal CPI_X_PC_INTERNAL_9 : std_logic ;
  signal CPI_X_PC_INTERNAL_10 : std_logic ;
  signal CPI_X_PC_INTERNAL_11 : std_logic ;
  signal CPI_X_PC_INTERNAL_12 : std_logic ;
  signal CPI_X_PC_INTERNAL_13 : std_logic ;
  signal CPI_X_PC_INTERNAL_14 : std_logic ;
  signal CPI_X_PC_INTERNAL_15 : std_logic ;
  signal CPI_X_PC_INTERNAL_16 : std_logic ;
  signal CPI_X_PC_INTERNAL_17 : std_logic ;
  signal CPI_X_PC_INTERNAL_18 : std_logic ;
  signal CPI_X_PC_INTERNAL_19 : std_logic ;
  signal CPI_X_PC_INTERNAL_20 : std_logic ;
  signal CPI_X_PC_INTERNAL_21 : std_logic ;
  signal CPI_X_PC_INTERNAL_22 : std_logic ;
  signal CPI_X_PC_INTERNAL_23 : std_logic ;
  signal CPI_X_PC_INTERNAL_24 : std_logic ;
  signal CPI_X_PC_INTERNAL_25 : std_logic ;
  signal CPI_X_PC_INTERNAL_26 : std_logic ;
  signal CPI_X_PC_INTERNAL_27 : std_logic ;
  signal CPI_X_PC_INTERNAL_28 : std_logic ;
  signal CPI_X_PC_INTERNAL_29 : std_logic ;
  signal CPI_X_PC_INTERNAL_30 : std_logic ;
  signal CPI_X_INST_INTERNAL : std_logic ;
  signal CPI_X_INST_INTERNAL_0 : std_logic ;
  signal CPI_X_INST_INTERNAL_1 : std_logic ;
  signal CPI_X_INST_INTERNAL_2 : std_logic ;
  signal CPI_X_INST_INTERNAL_3 : std_logic ;
  signal CPI_X_INST_INTERNAL_4 : std_logic ;
  signal CPI_X_INST_INTERNAL_5 : std_logic ;
  signal CPI_X_INST_INTERNAL_6 : std_logic ;
  signal CPI_X_INST_INTERNAL_7 : std_logic ;
  signal CPI_X_INST_INTERNAL_8 : std_logic ;
  signal CPI_X_INST_INTERNAL_9 : std_logic ;
  signal CPI_X_INST_INTERNAL_10 : std_logic ;
  signal CPI_X_INST_INTERNAL_11 : std_logic ;
  signal CPI_X_INST_INTERNAL_12 : std_logic ;
  signal CPI_X_INST_INTERNAL_13 : std_logic ;
  signal CPI_X_INST_INTERNAL_14 : std_logic ;
  signal CPI_X_INST_INTERNAL_15 : std_logic ;
  signal CPI_X_INST_INTERNAL_16 : std_logic ;
  signal CPI_X_INST_INTERNAL_17 : std_logic ;
  signal CPI_X_INST_INTERNAL_18 : std_logic ;
  signal CPI_X_INST_INTERNAL_19 : std_logic ;
  signal CPI_X_INST_INTERNAL_20 : std_logic ;
  signal CPI_X_INST_INTERNAL_21 : std_logic ;
  signal CPI_X_INST_INTERNAL_22 : std_logic ;
  signal CPI_X_INST_INTERNAL_23 : std_logic ;
  signal CPI_X_INST_INTERNAL_24 : std_logic ;
  signal CPI_X_INST_INTERNAL_25 : std_logic ;
  signal CPI_X_INST_INTERNAL_26 : std_logic ;
  signal CPI_X_INST_INTERNAL_27 : std_logic ;
  signal CPI_X_INST_INTERNAL_28 : std_logic ;
  signal CPI_X_INST_INTERNAL_29 : std_logic ;
  signal CPI_X_INST_INTERNAL_30 : std_logic ;
  signal CPI_X_CNT_INTERNAL : std_logic ;
  signal CPI_X_CNT_INTERNAL_0 : std_logic ;
  signal CPI_X_TRAP_INTERNAL : std_logic ;
  signal CPI_X_ANNUL_INTERNAL : std_logic ;
  signal CPI_X_PV_INTERNAL : std_logic ;
  signal CPI_LDDATA_INTERNAL : std_logic ;
  signal CPI_LDDATA_INTERNAL_0 : std_logic ;
  signal CPI_LDDATA_INTERNAL_1 : std_logic ;
  signal CPI_LDDATA_INTERNAL_2 : std_logic ;
  signal CPI_LDDATA_INTERNAL_3 : std_logic ;
  signal CPI_LDDATA_INTERNAL_4 : std_logic ;
  signal CPI_LDDATA_INTERNAL_5 : std_logic ;
  signal CPI_LDDATA_INTERNAL_6 : std_logic ;
  signal CPI_LDDATA_INTERNAL_7 : std_logic ;
  signal CPI_LDDATA_INTERNAL_8 : std_logic ;
  signal CPI_LDDATA_INTERNAL_9 : std_logic ;
  signal CPI_LDDATA_INTERNAL_10 : std_logic ;
  signal CPI_LDDATA_INTERNAL_11 : std_logic ;
  signal CPI_LDDATA_INTERNAL_12 : std_logic ;
  signal CPI_LDDATA_INTERNAL_13 : std_logic ;
  signal CPI_LDDATA_INTERNAL_14 : std_logic ;
  signal CPI_LDDATA_INTERNAL_15 : std_logic ;
  signal CPI_LDDATA_INTERNAL_16 : std_logic ;
  signal CPI_LDDATA_INTERNAL_17 : std_logic ;
  signal CPI_LDDATA_INTERNAL_18 : std_logic ;
  signal CPI_LDDATA_INTERNAL_19 : std_logic ;
  signal CPI_LDDATA_INTERNAL_20 : std_logic ;
  signal CPI_LDDATA_INTERNAL_21 : std_logic ;
  signal CPI_LDDATA_INTERNAL_22 : std_logic ;
  signal CPI_LDDATA_INTERNAL_23 : std_logic ;
  signal CPI_LDDATA_INTERNAL_24 : std_logic ;
  signal CPI_LDDATA_INTERNAL_25 : std_logic ;
  signal CPI_LDDATA_INTERNAL_26 : std_logic ;
  signal CPI_LDDATA_INTERNAL_27 : std_logic ;
  signal CPI_LDDATA_INTERNAL_28 : std_logic ;
  signal CPI_LDDATA_INTERNAL_29 : std_logic ;
  signal CPI_LDDATA_INTERNAL_30 : std_logic ;
  signal CPI_DBG_ENABLE_INTERNAL : std_logic ;
  signal CPI_DBG_WRITE_INTERNAL : std_logic ;
  signal CPI_DBG_FSR_INTERNAL : std_logic ;
  signal CPI_DBG_ADDR_INTERNAL : std_logic ;
  signal CPI_DBG_ADDR_INTERNAL_0 : std_logic ;
  signal CPI_DBG_ADDR_INTERNAL_1 : std_logic ;
  signal CPI_DBG_ADDR_INTERNAL_2 : std_logic ;
  signal CPI_DBG_ADDR_INTERNAL_3 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_0 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_1 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_2 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_3 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_4 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_5 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_6 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_7 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_8 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_9 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_10 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_11 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_12 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_13 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_14 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_15 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_16 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_17 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_18 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_19 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_20 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_21 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_22 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_23 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_24 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_25 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_26 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_27 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_28 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_29 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_30 : std_logic ;
  signal RFO1_DATA1_INTERNAL : std_logic ;
  signal RFO1_DATA1_INTERNAL_0 : std_logic ;
  signal RFO1_DATA1_INTERNAL_1 : std_logic ;
  signal RFO1_DATA1_INTERNAL_2 : std_logic ;
  signal RFO1_DATA1_INTERNAL_3 : std_logic ;
  signal RFO1_DATA1_INTERNAL_4 : std_logic ;
  signal RFO1_DATA1_INTERNAL_5 : std_logic ;
  signal RFO1_DATA1_INTERNAL_6 : std_logic ;
  signal RFO1_DATA1_INTERNAL_7 : std_logic ;
  signal RFO1_DATA1_INTERNAL_8 : std_logic ;
  signal RFO1_DATA1_INTERNAL_9 : std_logic ;
  signal RFO1_DATA1_INTERNAL_10 : std_logic ;
  signal RFO1_DATA1_INTERNAL_11 : std_logic ;
  signal RFO1_DATA1_INTERNAL_12 : std_logic ;
  signal RFO1_DATA1_INTERNAL_13 : std_logic ;
  signal RFO1_DATA1_INTERNAL_14 : std_logic ;
  signal RFO1_DATA1_INTERNAL_15 : std_logic ;
  signal RFO1_DATA1_INTERNAL_16 : std_logic ;
  signal RFO1_DATA1_INTERNAL_17 : std_logic ;
  signal RFO1_DATA1_INTERNAL_18 : std_logic ;
  signal RFO1_DATA1_INTERNAL_19 : std_logic ;
  signal RFO1_DATA1_INTERNAL_20 : std_logic ;
  signal RFO1_DATA1_INTERNAL_21 : std_logic ;
  signal RFO1_DATA1_INTERNAL_22 : std_logic ;
  signal RFO1_DATA1_INTERNAL_23 : std_logic ;
  signal RFO1_DATA1_INTERNAL_24 : std_logic ;
  signal RFO1_DATA1_INTERNAL_25 : std_logic ;
  signal RFO1_DATA1_INTERNAL_26 : std_logic ;
  signal RFO1_DATA1_INTERNAL_27 : std_logic ;
  signal RFO1_DATA1_INTERNAL_28 : std_logic ;
  signal RFO1_DATA1_INTERNAL_29 : std_logic ;
  signal RFO1_DATA1_INTERNAL_30 : std_logic ;
  signal RFO1_DATA2_INTERNAL : std_logic ;
  signal RFO1_DATA2_INTERNAL_0 : std_logic ;
  signal RFO1_DATA2_INTERNAL_1 : std_logic ;
  signal RFO1_DATA2_INTERNAL_2 : std_logic ;
  signal RFO1_DATA2_INTERNAL_3 : std_logic ;
  signal RFO1_DATA2_INTERNAL_4 : std_logic ;
  signal RFO1_DATA2_INTERNAL_5 : std_logic ;
  signal RFO1_DATA2_INTERNAL_6 : std_logic ;
  signal RFO1_DATA2_INTERNAL_7 : std_logic ;
  signal RFO1_DATA2_INTERNAL_8 : std_logic ;
  signal RFO1_DATA2_INTERNAL_9 : std_logic ;
  signal RFO1_DATA2_INTERNAL_10 : std_logic ;
  signal RFO1_DATA2_INTERNAL_11 : std_logic ;
  signal RFO1_DATA2_INTERNAL_12 : std_logic ;
  signal RFO1_DATA2_INTERNAL_13 : std_logic ;
  signal RFO1_DATA2_INTERNAL_14 : std_logic ;
  signal RFO1_DATA2_INTERNAL_15 : std_logic ;
  signal RFO1_DATA2_INTERNAL_16 : std_logic ;
  signal RFO1_DATA2_INTERNAL_17 : std_logic ;
  signal RFO1_DATA2_INTERNAL_18 : std_logic ;
  signal RFO1_DATA2_INTERNAL_19 : std_logic ;
  signal RFO1_DATA2_INTERNAL_20 : std_logic ;
  signal RFO1_DATA2_INTERNAL_21 : std_logic ;
  signal RFO1_DATA2_INTERNAL_22 : std_logic ;
  signal RFO1_DATA2_INTERNAL_23 : std_logic ;
  signal RFO1_DATA2_INTERNAL_24 : std_logic ;
  signal RFO1_DATA2_INTERNAL_25 : std_logic ;
  signal RFO1_DATA2_INTERNAL_26 : std_logic ;
  signal RFO1_DATA2_INTERNAL_27 : std_logic ;
  signal RFO1_DATA2_INTERNAL_28 : std_logic ;
  signal RFO1_DATA2_INTERNAL_29 : std_logic ;
  signal RFO1_DATA2_INTERNAL_30 : std_logic ;
  signal RFO2_DATA1_INTERNAL : std_logic ;
  signal RFO2_DATA1_INTERNAL_0 : std_logic ;
  signal RFO2_DATA1_INTERNAL_1 : std_logic ;
  signal RFO2_DATA1_INTERNAL_2 : std_logic ;
  signal RFO2_DATA1_INTERNAL_3 : std_logic ;
  signal RFO2_DATA1_INTERNAL_4 : std_logic ;
  signal RFO2_DATA1_INTERNAL_5 : std_logic ;
  signal RFO2_DATA1_INTERNAL_6 : std_logic ;
  signal RFO2_DATA1_INTERNAL_7 : std_logic ;
  signal RFO2_DATA1_INTERNAL_8 : std_logic ;
  signal RFO2_DATA1_INTERNAL_9 : std_logic ;
  signal RFO2_DATA1_INTERNAL_10 : std_logic ;
  signal RFO2_DATA1_INTERNAL_11 : std_logic ;
  signal RFO2_DATA1_INTERNAL_12 : std_logic ;
  signal RFO2_DATA1_INTERNAL_13 : std_logic ;
  signal RFO2_DATA1_INTERNAL_14 : std_logic ;
  signal RFO2_DATA1_INTERNAL_15 : std_logic ;
  signal RFO2_DATA1_INTERNAL_16 : std_logic ;
  signal RFO2_DATA1_INTERNAL_17 : std_logic ;
  signal RFO2_DATA1_INTERNAL_18 : std_logic ;
  signal RFO2_DATA1_INTERNAL_19 : std_logic ;
  signal RFO2_DATA1_INTERNAL_20 : std_logic ;
  signal RFO2_DATA1_INTERNAL_21 : std_logic ;
  signal RFO2_DATA1_INTERNAL_22 : std_logic ;
  signal RFO2_DATA1_INTERNAL_23 : std_logic ;
  signal RFO2_DATA1_INTERNAL_24 : std_logic ;
  signal RFO2_DATA1_INTERNAL_25 : std_logic ;
  signal RFO2_DATA1_INTERNAL_26 : std_logic ;
  signal RFO2_DATA1_INTERNAL_27 : std_logic ;
  signal RFO2_DATA1_INTERNAL_28 : std_logic ;
  signal RFO2_DATA1_INTERNAL_29 : std_logic ;
  signal RFO2_DATA1_INTERNAL_30 : std_logic ;
  signal RFO2_DATA2_INTERNAL : std_logic ;
  signal RFO2_DATA2_INTERNAL_0 : std_logic ;
  signal RFO2_DATA2_INTERNAL_1 : std_logic ;
  signal RFO2_DATA2_INTERNAL_2 : std_logic ;
  signal RFO2_DATA2_INTERNAL_3 : std_logic ;
  signal RFO2_DATA2_INTERNAL_4 : std_logic ;
  signal RFO2_DATA2_INTERNAL_5 : std_logic ;
  signal RFO2_DATA2_INTERNAL_6 : std_logic ;
  signal RFO2_DATA2_INTERNAL_7 : std_logic ;
  signal RFO2_DATA2_INTERNAL_8 : std_logic ;
  signal RFO2_DATA2_INTERNAL_9 : std_logic ;
  signal RFO2_DATA2_INTERNAL_10 : std_logic ;
  signal RFO2_DATA2_INTERNAL_11 : std_logic ;
  signal RFO2_DATA2_INTERNAL_12 : std_logic ;
  signal RFO2_DATA2_INTERNAL_13 : std_logic ;
  signal RFO2_DATA2_INTERNAL_14 : std_logic ;
  signal RFO2_DATA2_INTERNAL_15 : std_logic ;
  signal RFO2_DATA2_INTERNAL_16 : std_logic ;
  signal RFO2_DATA2_INTERNAL_17 : std_logic ;
  signal RFO2_DATA2_INTERNAL_18 : std_logic ;
  signal RFO2_DATA2_INTERNAL_19 : std_logic ;
  signal RFO2_DATA2_INTERNAL_20 : std_logic ;
  signal RFO2_DATA2_INTERNAL_21 : std_logic ;
  signal RFO2_DATA2_INTERNAL_22 : std_logic ;
  signal RFO2_DATA2_INTERNAL_23 : std_logic ;
  signal RFO2_DATA2_INTERNAL_24 : std_logic ;
  signal RFO2_DATA2_INTERNAL_25 : std_logic ;
  signal RFO2_DATA2_INTERNAL_26 : std_logic ;
  signal RFO2_DATA2_INTERNAL_27 : std_logic ;
  signal RFO2_DATA2_INTERNAL_28 : std_logic ;
  signal RFO2_DATA2_INTERNAL_29 : std_logic ;
  signal RFO2_DATA2_INTERNAL_30 : std_logic ;
  signal VCC : std_logic ;
  signal GND : std_logic ;
  signal \GRLFPC2_0.FPI.START\ : std_logic ;
  signal \GRLFPC2_0.FPI.RST\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\ : std_logic ;
  signal \GRLFPC2_0.R.I.EXEC\ : std_logic ;
  signal \GRLFPC2_0.R.X.LD\ : std_logic ;
  signal \GRLFPC2_0.R.X.AFSR\ : std_logic ;
  signal \GRLFPC2_0.R.X.SEQERR\ : std_logic ;
  signal \GRLFPC2_0.R.X.FPOP\ : std_logic ;
  signal \GRLFPC2_0.R.MK.HOLDN1\ : std_logic ;
  signal \GRLFPC2_0.R.E.FPOP\ : std_logic ;
  signal \GRLFPC2_0.R.M.FPOP\ : std_logic ;
  signal \GRLFPC2_0.R.MK.HOLDN2\ : std_logic ;
  signal \GRLFPC2_0.R.I.V\ : std_logic ;
  signal \GRLFPC2_0.R.M.LD\ : std_logic ;
  signal \GRLFPC2_0.R.E.LD\ : std_logic ;
  signal \GRLFPC2_0.R.A.LD\ : std_logic ;
  signal \GRLFPC2_0.R.A.FPOP\ : std_logic ;
  signal \GRLFPC2_0.R.X.AFQ\ : std_logic ;
  signal \GRLFPC2_0.R.I.RDD\ : std_logic ;
  signal \GRLFPC2_0.R.X.RDD\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.NONSTD\ : std_logic ;
  signal \GRLFPC2_0.COMB.RS2D_1\ : std_logic ;
  signal \GRLFPC2_0.N_554\ : std_logic ;
  signal \GRLFPC2_0.N_557\ : std_logic ;
  signal \GRLFPC2_0.N_558\ : std_logic ;
  signal \GRLFPC2_0.N_559\ : std_logic ;
  signal \GRLFPC2_0.N_95\ : std_logic ;
  signal \GRLFPC2_0.N_96\ : std_logic ;
  signal \GRLFPC2_0.N_97\ : std_logic ;
  signal \GRLFPC2_0.N_98\ : std_logic ;
  signal \GRLFPC2_0.N_99\ : std_logic ;
  signal \GRLFPC2_0.N_100\ : std_logic ;
  signal \GRLFPC2_0.N_101\ : std_logic ;
  signal \GRLFPC2_0.N_102\ : std_logic ;
  signal \GRLFPC2_0.N_103\ : std_logic ;
  signal \GRLFPC2_0.N_104\ : std_logic ;
  signal \GRLFPC2_0.N_105\ : std_logic ;
  signal \GRLFPC2_0.N_106\ : std_logic ;
  signal \GRLFPC2_0.N_107\ : std_logic ;
  signal \GRLFPC2_0.N_108\ : std_logic ;
  signal \GRLFPC2_0.N_109\ : std_logic ;
  signal \GRLFPC2_0.N_110\ : std_logic ;
  signal \GRLFPC2_0.N_111\ : std_logic ;
  signal \GRLFPC2_0.N_112\ : std_logic ;
  signal \GRLFPC2_0.N_113\ : std_logic ;
  signal \GRLFPC2_0.N_114\ : std_logic ;
  signal \GRLFPC2_0.N_115\ : std_logic ;
  signal \GRLFPC2_0.N_116\ : std_logic ;
  signal \GRLFPC2_0.N_117\ : std_logic ;
  signal \GRLFPC2_0.N_118\ : std_logic ;
  signal \GRLFPC2_0.N_119\ : std_logic ;
  signal \GRLFPC2_0.N_120\ : std_logic ;
  signal \GRLFPC2_0.N_121\ : std_logic ;
  signal \GRLFPC2_0.N_122\ : std_logic ;
  signal \GRLFPC2_0.N_123\ : std_logic ;
  signal \GRLFPC2_0.N_124\ : std_logic ;
  signal \GRLFPC2_0.N_125\ : std_logic ;
  signal \GRLFPC2_0.N_126\ : std_logic ;
  signal \GRLFPC2_0.N_127\ : std_logic ;
  signal \GRLFPC2_0.N_128\ : std_logic ;
  signal \GRLFPC2_0.N_129\ : std_logic ;
  signal \GRLFPC2_0.N_130\ : std_logic ;
  signal \GRLFPC2_0.N_131\ : std_logic ;
  signal \GRLFPC2_0.N_132\ : std_logic ;
  signal \GRLFPC2_0.N_133\ : std_logic ;
  signal \GRLFPC2_0.N_134\ : std_logic ;
  signal \GRLFPC2_0.N_135\ : std_logic ;
  signal \GRLFPC2_0.N_136\ : std_logic ;
  signal \GRLFPC2_0.N_137\ : std_logic ;
  signal \GRLFPC2_0.R.MK.RST\ : std_logic ;
  signal \GRLFPC2_0.COMB.ANNULFPU_1_O\ : std_logic ;
  signal \GRLFPC2_0.R.MK.HOLDN2_O\ : std_logic ;
  signal \GRLFPC2_0.R.MK.RST_O_0\ : std_logic ;
  signal \GRLFPC2_0.R.MK.RST2\ : std_logic ;
  signal \GRLFPC2_0.R.MK.RST2_O\ : std_logic ;
  signal \GRLFPC2_0.FPO.BUSY_O_0\ : std_logic ;
  signal \GRLFPC2_0.R.MK.HOLDN1_O_0\ : std_logic ;
  signal \GRLFPC2_0.R.MK.HOLDN2_O_0\ : std_logic ;
  signal \GRLFPC2_0.R.MK.RST2_O_0\ : std_logic ;
  signal \GRLFPC2_0.HOLDN_O\ : std_logic ;
  signal \GRLFPC2_0.COMB.LOCKGEN.LOCKI_O_3\ : std_logic ;
  signal \GRLFPC2_0.R.MK.BUSY_O\ : std_logic ;
  signal \GRLFPC2_0.COMB.LOCKGEN.LOCKI_O\ : std_logic ;
  signal \GRLFPC2_0.COMB.ANNULFPU_1_O_0\ : std_logic ;
  signal \GRLFPC2_0.N_835\ : std_logic ;
  signal \GRLFPC2_0.COMB.FPDECODE.ST_O\ : std_logic ;
  signal \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\ : std_logic ;
  signal \GRLFPC2_0.R.A.AFSR_O\ : std_logic ;
  signal \GRLFPC2_0.N_553\ : std_logic ;
  signal \GRLFPC2_0.N_1837_O\ : std_logic ;
  signal \GRLFPC2_0.R.A.RS1D\ : std_logic ;
  signal \GRLFPC2_0.R.A.RS2D\ : std_logic ;
  signal \GRLFPC2_0.R.A.AFQ_O\ : std_logic ;
  signal \GRLFPC2_0.R.E.AFSR_O\ : std_logic ;
  signal \GRLFPC2_0.R.E.AFQ_O\ : std_logic ;
  signal \GRLFPC2_0.N_1829_O\ : std_logic ;
  signal \GRLFPC2_0.N_1105\ : std_logic ;
  signal \GRLFPC2_0.N_1000\ : std_logic ;
  signal \GRLFPC2_0.N_2101\ : std_logic ;
  signal \GRLFPC2_0.N_2111\ : std_logic ;
  signal \GRLFPC2_0.N_2115\ : std_logic ;
  signal \GRLFPC2_0.COMB.ANNULFPU_1\ : std_logic ;
  signal \GRLFPC2_0.COMB.RS1D_1\ : std_logic ;
  signal \GRLFPC2_0.N_884\ : std_logic ;
  signal \GRLFPC2_0.N_620\ : std_logic ;
  signal \GRLFPC2_0.N_925\ : std_logic ;
  signal \GRLFPC2_0.N_889\ : std_logic ;
  signal \GRLFPC2_0.N_178\ : std_logic ;
  signal \GRLFPC2_0.N_3418\ : std_logic ;
  signal \GRLFPC2_0.N_92\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5410\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5391\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN25_NOTPROP\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_954\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4459\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7248\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7259\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7260\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7272\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7274\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10026\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10027\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10028\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10029\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10030\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10031\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10032\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10033\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10034\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10035\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10036\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10037\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10038\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10039\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10040\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10041\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10042\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10043\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10044\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10045\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10046\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10047\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10048\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10049\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10050\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10051\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10052\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10053\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10054\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10055\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10056\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10057\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10058\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10059\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10060\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10061\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10062\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10063\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10064\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10065\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10066\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10067\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10068\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10069\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10070\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10071\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10072\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10073\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10074\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10076\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10077\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10078\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10079\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10080\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10081\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10082\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10085\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10086\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10087\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10088\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10089\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10090\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10091\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10092\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10093\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10094\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10095\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10096\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10097\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10098\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10099\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10100\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10101\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10102\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10103\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10104\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10105\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10106\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10107\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10108\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10109\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10110\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10111\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10112\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10113\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10114\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10115\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10116\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10117\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10118\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10119\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10120\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10121\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10122\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10123\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10124\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10125\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10126\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10127\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10128\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10129\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10130\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10131\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10132\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10133\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10134\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10135\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10136\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10137\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10138\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10139\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10140\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10141\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10142\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10560\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_I\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3926\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.TEMP\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_377\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2765\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2807\ : std_logic ;
  signal N_1 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1780_I\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.UN36_PCTRL_NEW_I\ : std_logic ;
  signal N_26534 : std_logic ;
  signal N_26535 : std_logic ;
  signal N_26536 : std_logic ;
  signal N_26537 : std_logic ;
  signal N_26538 : std_logic ;
  signal N_26539 : std_logic ;
  signal N_26540 : std_logic ;
  signal N_26541 : std_logic ;
  signal N_26542 : std_logic ;
  signal N_26543 : std_logic ;
  signal N_26544 : std_logic ;
  signal N_26545 : std_logic ;
  signal N_26546 : std_logic ;
  signal N_26547 : std_logic ;
  signal N_26548 : std_logic ;
  signal N_26549 : std_logic ;
  signal N_26550 : std_logic ;
  signal N_26551 : std_logic ;
  signal N_26552 : std_logic ;
  signal N_26553 : std_logic ;
  signal N_26554 : std_logic ;
  signal N_26555 : std_logic ;
  signal N_26556 : std_logic ;
  signal N_26557 : std_logic ;
  signal N_26558 : std_logic ;
  signal N_26559 : std_logic ;
  signal N_26560 : std_logic ;
  signal N_26561 : std_logic ;
  signal N_26562 : std_logic ;
  signal N_26563 : std_logic ;
  signal N_26564 : std_logic ;
  signal N_26565 : std_logic ;
  signal N_26566 : std_logic ;
  signal N_26567 : std_logic ;
  signal N_26568 : std_logic ;
  signal N_26569 : std_logic ;
  signal N_26570 : std_logic ;
  signal N_26571 : std_logic ;
  signal N_26572 : std_logic ;
  signal N_26573 : std_logic ;
  signal N_26574 : std_logic ;
  signal N_26575 : std_logic ;
  signal N_26576 : std_logic ;
  signal N_26577 : std_logic ;
  signal N_26578 : std_logic ;
  signal N_26579 : std_logic ;
  signal N_26580 : std_logic ;
  signal N_26581 : std_logic ;
  signal N_26582 : std_logic ;
  signal N_26583 : std_logic ;
  signal N_26584 : std_logic ;
  signal N_26585 : std_logic ;
  signal N_26586 : std_logic ;
  signal N_26587 : std_logic ;
  signal N_26588 : std_logic ;
  signal N_26589 : std_logic ;
  signal N_26590 : std_logic ;
  signal N_26591 : std_logic ;
  signal N_26592 : std_logic ;
  signal N_28672 : std_logic ;
  signal N_28673 : std_logic ;
  signal N_28675 : std_logic ;
  signal N_28676 : std_logic ;
  signal N_28678 : std_logic ;
  signal N_28679 : std_logic ;
  signal N_28681 : std_logic ;
  signal N_28682 : std_logic ;
  signal N_28684 : std_logic ;
  signal N_28685 : std_logic ;
  signal N_28687 : std_logic ;
  signal N_28688 : std_logic ;
  signal N_28690 : std_logic ;
  signal N_28691 : std_logic ;
  signal N_28693 : std_logic ;
  signal N_28694 : std_logic ;
  signal N_28696 : std_logic ;
  signal N_28697 : std_logic ;
  signal N_28699 : std_logic ;
  signal N_28700 : std_logic ;
  signal N_28702 : std_logic ;
  signal N_28703 : std_logic ;
  signal N_28705 : std_logic ;
  signal N_28706 : std_logic ;
  signal N_28708 : std_logic ;
  signal N_28709 : std_logic ;
  signal N_28711 : std_logic ;
  signal N_28712 : std_logic ;
  signal N_28714 : std_logic ;
  signal N_28715 : std_logic ;
  signal N_28717 : std_logic ;
  signal N_28718 : std_logic ;
  signal N_28720 : std_logic ;
  signal N_28721 : std_logic ;
  signal N_28723 : std_logic ;
  signal N_28724 : std_logic ;
  signal N_28726 : std_logic ;
  signal N_28727 : std_logic ;
  signal N_28729 : std_logic ;
  signal N_28730 : std_logic ;
  signal N_28732 : std_logic ;
  signal N_28733 : std_logic ;
  signal N_28735 : std_logic ;
  signal N_28736 : std_logic ;
  signal N_28738 : std_logic ;
  signal N_28739 : std_logic ;
  signal N_28741 : std_logic ;
  signal N_28742 : std_logic ;
  signal N_28744 : std_logic ;
  signal N_28745 : std_logic ;
  signal N_28747 : std_logic ;
  signal N_28748 : std_logic ;
  signal N_28750 : std_logic ;
  signal N_28751 : std_logic ;
  signal N_28753 : std_logic ;
  signal N_28754 : std_logic ;
  signal N_28756 : std_logic ;
  signal N_28757 : std_logic ;
  signal N_28759 : std_logic ;
  signal N_28760 : std_logic ;
  signal N_28762 : std_logic ;
  signal N_28763 : std_logic ;
  signal N_28765 : std_logic ;
  signal N_28766 : std_logic ;
  signal N_28768 : std_logic ;
  signal N_28769 : std_logic ;
  signal N_28771 : std_logic ;
  signal N_28772 : std_logic ;
  signal N_28774 : std_logic ;
  signal N_28775 : std_logic ;
  signal N_28777 : std_logic ;
  signal N_28778 : std_logic ;
  signal N_28780 : std_logic ;
  signal N_28781 : std_logic ;
  signal N_28783 : std_logic ;
  signal N_28784 : std_logic ;
  signal N_28786 : std_logic ;
  signal N_28787 : std_logic ;
  signal N_28789 : std_logic ;
  signal N_28790 : std_logic ;
  signal N_28792 : std_logic ;
  signal N_28793 : std_logic ;
  signal N_28795 : std_logic ;
  signal N_28796 : std_logic ;
  signal N_28798 : std_logic ;
  signal N_28799 : std_logic ;
  signal N_28801 : std_logic ;
  signal N_28802 : std_logic ;
  signal N_28804 : std_logic ;
  signal N_28805 : std_logic ;
  signal N_28807 : std_logic ;
  signal N_28808 : std_logic ;
  signal N_28810 : std_logic ;
  signal N_28811 : std_logic ;
  signal N_28813 : std_logic ;
  signal N_28814 : std_logic ;
  signal N_28816 : std_logic ;
  signal N_28817 : std_logic ;
  signal N_28819 : std_logic ;
  signal N_28820 : std_logic ;
  signal N_28822 : std_logic ;
  signal N_28823 : std_logic ;
  signal N_28825 : std_logic ;
  signal N_28826 : std_logic ;
  signal N_28828 : std_logic ;
  signal N_28829 : std_logic ;
  signal N_28831 : std_logic ;
  signal N_28832 : std_logic ;
  signal N_28834 : std_logic ;
  signal N_28835 : std_logic ;
  signal N_28837 : std_logic ;
  signal N_28838 : std_logic ;
  signal N_28840 : std_logic ;
  signal N_28841 : std_logic ;
  signal N_28843 : std_logic ;
  signal N_28844 : std_logic ;
  signal N_28846 : std_logic ;
  signal N_28847 : std_logic ;
  signal N_28849 : std_logic ;
  signal N_28850 : std_logic ;
  signal N_28852 : std_logic ;
  signal N_28853 : std_logic ;
  signal N_28855 : std_logic ;
  signal N_28856 : std_logic ;
  signal N_28858 : std_logic ;
  signal N_28859 : std_logic ;
  signal N_28861 : std_logic ;
  signal N_28862 : std_logic ;
  signal N_28864 : std_logic ;
  signal N_28865 : std_logic ;
  signal N_28867 : std_logic ;
  signal N_28868 : std_logic ;
  signal N_28870 : std_logic ;
  signal N_28871 : std_logic ;
  signal N_28873 : std_logic ;
  signal N_28874 : std_logic ;
  signal N_28876 : std_logic ;
  signal N_28877 : std_logic ;
  signal N_28879 : std_logic ;
  signal N_28880 : std_logic ;
  signal N_28882 : std_logic ;
  signal N_28883 : std_logic ;
  signal N_28885 : std_logic ;
  signal N_28886 : std_logic ;
  signal N_28888 : std_logic ;
  signal N_28889 : std_logic ;
  signal N_28891 : std_logic ;
  signal N_28892 : std_logic ;
  signal N_28894 : std_logic ;
  signal N_28895 : std_logic ;
  signal N_28897 : std_logic ;
  signal N_28898 : std_logic ;
  signal N_28900 : std_logic ;
  signal N_28901 : std_logic ;
  signal N_28903 : std_logic ;
  signal N_28904 : std_logic ;
  signal N_28906 : std_logic ;
  signal N_28907 : std_logic ;
  signal N_28909 : std_logic ;
  signal N_28910 : std_logic ;
  signal N_28912 : std_logic ;
  signal N_28913 : std_logic ;
  signal N_28915 : std_logic ;
  signal N_28916 : std_logic ;
  signal N_28918 : std_logic ;
  signal N_28919 : std_logic ;
  signal N_28921 : std_logic ;
  signal N_28922 : std_logic ;
  signal N_28924 : std_logic ;
  signal N_28925 : std_logic ;
  signal N_28927 : std_logic ;
  signal N_28928 : std_logic ;
  signal N_28930 : std_logic ;
  signal N_28931 : std_logic ;
  signal N_28933 : std_logic ;
  signal N_28934 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2466_1\ : std_logic ;
  signal \GRLFPC2_0.R.MK.BUSY_4\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.I.EXEC_1_3\ : std_logic ;
  signal \GRLFPC2_0.N_50_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_47__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_44__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_43__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_41__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_40__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_39__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_35__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_30__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_24__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_23__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_22__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_21__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_20__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_16__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_15__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_14__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_8__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_2__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_1__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_372__G1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_319__G1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_318__G1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_317__G1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_316__G1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_258__N_5_I\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_176__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_175__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_57__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_54__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_53__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_52__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_51__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_50__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_49__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_48__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_47__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_46__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_45__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_44__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_43__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_42__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_41__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_40__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_39__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_38__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_37__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_36__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_35__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_34__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_33__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_32__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_31__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_30__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_29__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_28__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_27__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_26__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_25__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_24__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_23__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_22__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_21__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_20__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_19__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_18__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_17__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_16__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_15__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_14__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_13__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_11__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_10__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_9__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_8__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_7__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_6__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_5__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_4__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_3__G2\ : std_logic ;
  signal \GRLFPC2_0.R.M.AFQ_RET_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.M.AFSR_RET_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.COMB.FPDECODE.ST\ : std_logic ;
  signal \GRLFPC2_0.R.E.SEQERR_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.V.I.EXEC_0_SQMUXA\ : std_logic ;
  signal \GRLFPC2_0.R.A.RDD_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.A.LD_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.FTT_0_0_0__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.NONSTD_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.I.RDD_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.X.LD_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.X.FPOP_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.X.AFSR_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.X.AFQ_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.M.LD_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.M.FPOP_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.LD_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.E.FPOP_1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_0__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_1__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_2__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_3__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_4__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_5__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_6__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_7__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_8__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_9__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_10__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_11__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_12__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_13__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_14__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_15__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_16__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_17__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_18__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_19__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_20__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_21__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_22__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_23__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_24__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_25__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_26__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_27__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_28__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_29__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_30__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_31__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.RD_0_0_0__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.RD_0_0_1__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.TEM_1_0_0__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.TEM_1_0_1__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.TEM_1_0_2__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.TEM_1_0_3__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.TEM_1_0_4__G1\ : std_logic ;
  signal \GRLFPC2_0.R.STATE_0_0_0__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.FCC_0_0_0__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.FCC_0_0_1__G1\ : std_logic ;
  signal \GRLFPC2_0.R.I.CC_0_0_0__G2\ : std_logic ;
  signal \GRLFPC2_0.R.I.CC_0_0_1__G2\ : std_logic ;
  signal \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\ : std_logic ;
  signal \GRLFPC2_0.R.I.EXC_2_0_1__G2\ : std_logic ;
  signal \GRLFPC2_0.R.I.EXC_2_0_2__G2\ : std_logic ;
  signal \GRLFPC2_0.R.I.EXC_2_0_3__G2\ : std_logic ;
  signal \GRLFPC2_0.R.I.EXC_2_0_4__G2\ : std_logic ;
  signal N_35958 : std_logic ;
  signal N_35959 : std_logic ;
  signal N_36149 : std_logic ;
  signal N_36176 : std_logic ;
  signal N_36203 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6_I\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_48__I0_I_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__I0_I_0\ : std_logic ;
  signal N_36366 : std_logic ;
  signal N_36367 : std_logic ;
  signal N_36368 : std_logic ;
  signal N_36369 : std_logic ;
  signal N_36370 : std_logic ;
  signal N_36371 : std_logic ;
  signal N_36372 : std_logic ;
  signal N_36373 : std_logic ;
  signal N_36374 : std_logic ;
  signal N_36375 : std_logic ;
  signal \GRLFPC2_0.R.STATE_0_0_1__I0_I_1\ : std_logic ;
  signal N_36379 : std_logic ;
  signal N_36380 : std_logic ;
  signal N_36381 : std_logic ;
  signal N_36382 : std_logic ;
  signal \GRLFPC2_0.R.FSR.AEXC_1_0_0__I0_I_0\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.AEXC_1_0_1__I0_I_1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.AEXC_1_0_2__I0_I_0\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.AEXC_1_0_3__I0_I_1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.AEXC_1_0_4__I0_I_0\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.CEXC_1_0_0__I0_I_1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.CEXC_1_0_1__I0_I_0\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.CEXC_1_0_2__I0_I_1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.CEXC_1_0_3__I0_I_0\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.CEXC_1_0_4__I0_I_1\ : std_logic ;
  signal RST_INTERNAL : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\ : std_logic ;
  signal N_48774 : std_logic ;
  signal N_48775 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5330\ : std_logic ;
  signal \GRLFPC2_0.N_1093\ : std_logic ;
  signal \GRLFPC2_0.COMB.FPDECODE.RS1D5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5065\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5088\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN14_EXMIPTRLSBS\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M\ : std_logic ;
  signal N_31688 : std_logic ;
  signal N_31788 : std_logic ;
  signal N_33138_1 : std_logic ;
  signal N_32400 : std_logic ;
  signal N_32404 : std_logic ;
  signal N_32405 : std_logic ;
  signal N_32394_I : std_logic ;
  signal N_31919 : std_logic ;
  signal N_31944 : std_logic ;
  signal N_32426 : std_logic ;
  signal N_32428 : std_logic ;
  signal N_32434 : std_logic ;
  signal N_32425 : std_logic ;
  signal N_31810 : std_logic ;
  signal N_31766_1 : std_logic ;
  signal N_32120_1 : std_logic ;
  signal N_31811_2 : std_logic ;
  signal N_32136_1 : std_logic ;
  signal N_31813_2 : std_logic ;
  signal N_32340_1 : std_logic ;
  signal N_31766_2 : std_logic ;
  signal N_33063_1 : std_logic ;
  signal N_31919_1 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_320\ : std_logic ;
  signal N_31839_1 : std_logic ;
  signal N_31892 : std_logic ;
  signal N_32487_2 : std_logic ;
  signal N_27553_1 : std_logic ;
  signal N_32070_1 : std_logic ;
  signal N_32688_1 : std_logic ;
  signal N_32413_2 : std_logic ;
  signal N_32908_1 : std_logic ;
  signal N_32272_2 : std_logic ;
  signal N_32418_1 : std_logic ;
  signal N_32425_1 : std_logic ;
  signal N_32047_1 : std_logic ;
  signal N_31989_1 : std_logic ;
  signal N_31819_2 : std_logic ;
  signal N_32432 : std_logic ;
  signal N_32048_1 : std_logic ;
  signal N_32066_2 : std_logic ;
  signal N_32434_2 : std_logic ;
  signal N_32131_1 : std_logic ;
  signal N_32435_1 : std_logic ;
  signal N_32438_1 : std_logic ;
  signal N_32140_1 : std_logic ;
  signal N_33298 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2599\ : std_logic ;
  signal N_32673_I : std_logic ;
  signal N_32739 : std_logic ;
  signal N_28580_1 : std_logic ;
  signal N_31763_1 : std_logic ;
  signal N_33176 : std_logic ;
  signal N_31931 : std_logic ;
  signal N_31921 : std_logic ;
  signal N_32838 : std_logic ;
  signal N_32836 : std_logic ;
  signal N_32852 : std_logic ;
  signal N_32700 : std_logic ;
  signal N_32708 : std_logic ;
  signal N_32693 : std_logic ;
  signal N_31769_1 : std_logic ;
  signal N_31931_1 : std_logic ;
  signal N_32136_2 : std_logic ;
  signal N_31940_1 : std_logic ;
  signal N_32500_2 : std_logic ;
  signal N_32290_1 : std_logic ;
  signal N_32566_1 : std_logic ;
  signal N_31774_1 : std_logic ;
  signal N_33145_4 : std_logic ;
  signal N_32662_I : std_logic ;
  signal N_32220_1 : std_logic ;
  signal N_31723_1 : std_logic ;
  signal N_31718_1 : std_logic ;
  signal N_31765_1 : std_logic ;
  signal N_32712_3 : std_logic ;
  signal N_32064_1 : std_logic ;
  signal N_27297_1 : std_logic ;
  signal N_32839_3 : std_logic ;
  signal N_32841_2 : std_logic ;
  signal N_31808_1 : std_logic ;
  signal N_32848 : std_logic ;
  signal N_32069_2 : std_logic ;
  signal N_32632_1 : std_logic ;
  signal N_31886_2 : std_logic ;
  signal \GRLFPC2_0.N_1092\ : std_logic ;
  signal N_36334 : std_logic ;
  signal \GRLFPC2_0.N_896\ : std_logic ;
  signal \GRLFPC2_0.N_889_1\ : std_logic ;
  signal N_36289 : std_logic ;
  signal \GRLFPC2_0.N_93\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10906\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10909\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10913\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10916\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10918\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10920\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10924\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10927\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916\ : std_logic ;
  signal N_28949 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SFTLFT.AREGXORBREG_I_M\ : std_logic ;
  signal N_28946 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642\ : std_logic ;
  signal N_28950 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2555\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2645\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2477\ : std_logic ;
  signal \GRLFPC2_0.N_37\ : std_logic ;
  signal N_31775_1 : std_logic ;
  signal N_32894 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2706\ : std_logic ;
  signal N_32246 : std_logic ;
  signal N_32327 : std_logic ;
  signal \GRLFPC2_0.N_73\ : std_logic ;
  signal N_33352 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1941\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_596\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2359\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_523\ : std_logic ;
  signal N_31862 : std_logic ;
  signal N_32143 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1931\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1071\ : std_logic ;
  signal N_31762 : std_logic ;
  signal N_32483 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2407\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1937\ : std_logic ;
  signal N_32853 : std_logic ;
  signal N_32695 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3924\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9471\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1788\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2659\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2582_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2622_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2560\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2674\ : std_logic ;
  signal N_27776_2 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2321\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2796\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2319\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2318\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2576_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_247\ : std_logic ;
  signal N_28030_I : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1958\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1956\ : std_logic ;
  signal N_31715_1 : std_logic ;
  signal N_31713 : std_logic ;
  signal N_31714 : std_logic ;
  signal N_31753 : std_logic ;
  signal N_31922 : std_logic ;
  signal N_31768_1 : std_logic ;
  signal N_31991 : std_logic ;
  signal N_32050 : std_logic ;
  signal N_32645_3 : std_logic ;
  signal N_32050_1 : std_logic ;
  signal N_32128_1 : std_logic ;
  signal N_32134_2 : std_logic ;
  signal N_32198_1 : std_logic ;
  signal N_32232 : std_logic ;
  signal N_32210 : std_logic ;
  signal N_32273 : std_logic ;
  signal N_31819_1 : std_logic ;
  signal N_32712_1 : std_logic ;
  signal N_32275 : std_logic ;
  signal N_32124_2 : std_logic ;
  signal N_32345 : std_logic ;
  signal N_33057_1 : std_logic ;
  signal N_32345_2 : std_logic ;
  signal N_32436 : std_logic ;
  signal N_32485 : std_logic ;
  signal N_31999_1 : std_logic ;
  signal N_32485_1 : std_logic ;
  signal N_31838_1 : std_logic ;
  signal N_32773 : std_logic ;
  signal N_31996_1 : std_logic ;
  signal N_32901 : std_logic ;
  signal N_32903 : std_logic ;
  signal N_31762_1 : std_logic ;
  signal N_32983 : std_logic ;
  signal N_32984 : std_logic ;
  signal N_32985 : std_logic ;
  signal N_32705_1 : std_logic ;
  signal N_32142_1 : std_logic ;
  signal N_33058 : std_logic ;
  signal N_33129 : std_logic ;
  signal N_33131 : std_logic ;
  signal N_28591_1 : std_logic ;
  signal N_33255 : std_logic ;
  signal N_33232 : std_logic ;
  signal N_33256 : std_logic ;
  signal N_31865_1 : std_logic ;
  signal N_33367 : std_logic ;
  signal N_31941_1 : std_logic ;
  signal N_32344_1 : std_logic ;
  signal N_33360 : std_logic ;
  signal N_33359 : std_logic ;
  signal N_33372 : std_logic ;
  signal N_33357 : std_logic ;
  signal N_33356 : std_logic ;
  signal N_33136_2 : std_logic ;
  signal N_31718_2 : std_logic ;
  signal N_33355 : std_logic ;
  signal N_31864_1 : std_logic ;
  signal N_33333 : std_logic ;
  signal N_32230 : std_logic ;
  signal N_32786_1 : std_logic ;
  signal N_33316 : std_logic ;
  signal N_33314_4 : std_logic ;
  signal N_27929_1 : std_logic ;
  signal N_32093 : std_logic ;
  signal N_33312 : std_logic ;
  signal N_33312_2 : std_logic ;
  signal N_33311 : std_logic ;
  signal N_33310 : std_logic ;
  signal N_33277 : std_logic ;
  signal N_33276 : std_logic ;
  signal N_33275 : std_logic ;
  signal N_33275_1 : std_logic ;
  signal N_33274 : std_logic ;
  signal N_33076_1 : std_logic ;
  signal N_33271 : std_logic ;
  signal N_33268 : std_logic ;
  signal N_32619_1 : std_logic ;
  signal N_33264_2 : std_logic ;
  signal N_33261 : std_logic ;
  signal N_33260 : std_logic ;
  signal N_27758_I : std_logic ;
  signal N_33259 : std_logic ;
  signal N_32885_I : std_logic ;
  signal N_32708_2 : std_logic ;
  signal N_33209 : std_logic ;
  signal N_33208 : std_logic ;
  signal N_32278_2 : std_logic ;
  signal N_33207_1 : std_logic ;
  signal N_33206 : std_logic ;
  signal N_33136_1 : std_logic ;
  signal N_33203 : std_logic ;
  signal N_33202 : std_logic ;
  signal N_32422_1 : std_logic ;
  signal N_32530_I : std_logic ;
  signal N_33201 : std_logic ;
  signal N_32620_1 : std_logic ;
  signal N_33200 : std_logic ;
  signal N_33198 : std_logic ;
  signal N_33197 : std_logic ;
  signal N_33196 : std_logic ;
  signal N_32550_1 : std_logic ;
  signal N_33193 : std_logic ;
  signal N_31724_1 : std_logic ;
  signal N_33148 : std_logic ;
  signal N_33167 : std_logic ;
  signal N_33145 : std_logic ;
  signal N_33144 : std_logic ;
  signal N_33143 : std_logic ;
  signal N_33143_1 : std_logic ;
  signal N_33141_2 : std_logic ;
  signal N_33140 : std_logic ;
  signal N_33136 : std_logic ;
  signal N_33135 : std_logic ;
  signal N_33134_1 : std_logic ;
  signal N_33130 : std_logic ;
  signal N_32343_1 : std_logic ;
  signal N_33128 : std_logic ;
  signal N_33127 : std_logic ;
  signal N_32645_2 : std_logic ;
  signal N_33126 : std_logic ;
  signal N_33032 : std_logic ;
  signal N_33080 : std_logic ;
  signal N_33075 : std_logic ;
  signal N_33072 : std_logic ;
  signal N_32015_1 : std_logic ;
  signal N_33071_1 : std_logic ;
  signal N_33067 : std_logic ;
  signal N_33064 : std_logic ;
  signal N_33064_1 : std_logic ;
  signal N_33060 : std_logic ;
  signal N_33040 : std_logic ;
  signal N_33001_1 : std_logic ;
  signal N_33023 : std_logic ;
  signal N_32999 : std_logic ;
  signal N_32998 : std_logic ;
  signal N_32203_1 : std_logic ;
  signal N_32995_1 : std_logic ;
  signal N_32994 : std_logic ;
  signal N_32992 : std_logic ;
  signal N_32991 : std_logic ;
  signal N_31899_I : std_logic ;
  signal N_32986 : std_logic ;
  signal N_32980 : std_logic ;
  signal N_32932 : std_logic ;
  signal N_32925_2 : std_logic ;
  signal N_32922 : std_logic ;
  signal N_32914 : std_logic ;
  signal N_32913 : std_logic ;
  signal N_32912 : std_logic ;
  signal N_32911 : std_logic ;
  signal N_32909 : std_logic ;
  signal N_32908 : std_logic ;
  signal N_32907 : std_logic ;
  signal N_32906 : std_logic ;
  signal N_32905 : std_logic ;
  signal N_32904 : std_logic ;
  signal N_32849 : std_logic ;
  signal N_32846 : std_logic ;
  signal N_32841 : std_logic ;
  signal N_32840_3 : std_logic ;
  signal N_31691_I : std_logic ;
  signal N_32765 : std_logic ;
  signal N_32785 : std_logic ;
  signal N_32785_2 : std_logic ;
  signal N_32784 : std_logic ;
  signal N_32784_2 : std_logic ;
  signal N_32777 : std_logic ;
  signal N_32775 : std_logic ;
  signal N_32775_1 : std_logic ;
  signal N_32770 : std_logic ;
  signal N_32768 : std_logic ;
  signal N_32766 : std_logic ;
  signal N_32710 : std_logic ;
  signal N_32702 : std_logic ;
  signal N_32699 : std_logic ;
  signal N_32698 : std_logic ;
  signal N_31767_2 : std_logic ;
  signal N_32691 : std_logic ;
  signal N_32688 : std_logic ;
  signal N_32032_I : std_logic ;
  signal N_32641 : std_logic ;
  signal N_32628 : std_logic ;
  signal N_32627_1 : std_logic ;
  signal N_32626 : std_logic ;
  signal N_32625 : std_logic ;
  signal N_32624 : std_logic ;
  signal N_32622 : std_logic ;
  signal N_32621 : std_logic ;
  signal N_32620 : std_logic ;
  signal N_32587 : std_logic ;
  signal N_32586 : std_logic ;
  signal N_32567_2 : std_logic ;
  signal N_32564 : std_logic ;
  signal N_32563_2 : std_logic ;
  signal N_32559 : std_logic ;
  signal N_32558 : std_logic ;
  signal N_32553 : std_logic ;
  signal N_32552 : std_logic ;
  signal N_32551 : std_logic ;
  signal N_32549 : std_logic ;
  signal N_32548 : std_logic ;
  signal N_32546 : std_logic ;
  signal N_32545 : std_logic ;
  signal N_32500 : std_logic ;
  signal N_32498_4 : std_logic ;
  signal N_32497 : std_logic ;
  signal N_32496 : std_logic ;
  signal N_32492 : std_logic ;
  signal N_32487 : std_logic ;
  signal N_32484 : std_logic ;
  signal N_32427 : std_logic ;
  signal N_32424 : std_logic ;
  signal N_32423 : std_logic ;
  signal N_32390_I : std_logic ;
  signal N_32422 : std_logic ;
  signal N_32421 : std_logic ;
  signal N_32416 : std_logic ;
  signal N_32357 : std_logic ;
  signal N_32354 : std_logic ;
  signal N_32350 : std_logic ;
  signal N_32322_I : std_logic ;
  signal N_32348 : std_logic ;
  signal N_32347 : std_logic ;
  signal N_32346 : std_logic ;
  signal N_32343 : std_logic ;
  signal N_32341 : std_logic ;
  signal N_32340 : std_logic ;
  signal N_32336 : std_logic ;
  signal N_32289_2 : std_logic ;
  signal N_32287 : std_logic ;
  signal N_32281 : std_logic ;
  signal N_32280 : std_logic ;
  signal N_32279 : std_logic ;
  signal N_32279_3 : std_logic ;
  signal N_32277 : std_logic ;
  signal N_32274 : std_logic ;
  signal N_32272 : std_logic ;
  signal N_32221_1 : std_logic ;
  signal N_32217_1 : std_logic ;
  signal N_32209 : std_logic ;
  signal N_32207_1 : std_logic ;
  signal N_32206_2 : std_logic ;
  signal N_32200 : std_logic ;
  signal N_32199 : std_logic ;
  signal N_32197 : std_logic ;
  signal N_32196 : std_logic ;
  signal N_32195 : std_logic ;
  signal N_32194 : std_logic ;
  signal N_32141 : std_logic ;
  signal N_32139 : std_logic ;
  signal N_32136 : std_logic ;
  signal N_32135_2 : std_logic ;
  signal N_32133 : std_logic ;
  signal N_32131 : std_logic ;
  signal N_32130 : std_logic ;
  signal N_32127 : std_logic ;
  signal N_32126 : std_logic ;
  signal N_32124 : std_logic ;
  signal N_32122 : std_logic ;
  signal N_32120 : std_logic ;
  signal N_32064 : std_logic ;
  signal N_32061 : std_logic ;
  signal N_32020 : std_logic ;
  signal N_32057_2 : std_logic ;
  signal N_32056 : std_logic ;
  signal N_32022_I : std_logic ;
  signal N_32023 : std_logic ;
  signal N_32052 : std_logic ;
  signal N_32049 : std_logic ;
  signal N_32048 : std_logic ;
  signal N_32046 : std_logic ;
  signal N_31998 : std_logic ;
  signal N_31997 : std_logic ;
  signal N_31993 : std_logic ;
  signal N_31989 : std_logic ;
  signal N_31983 : std_logic ;
  signal N_31946 : std_logic ;
  signal N_31945 : std_logic ;
  signal N_31929 : std_logic ;
  signal N_31926 : std_logic ;
  signal N_31918 : std_logic ;
  signal N_31875 : std_logic ;
  signal N_31867 : std_logic ;
  signal N_31865 : std_logic ;
  signal N_31864 : std_logic ;
  signal N_31819 : std_logic ;
  signal N_31818 : std_logic ;
  signal N_31817 : std_logic ;
  signal N_31816_1 : std_logic ;
  signal N_31814 : std_logic ;
  signal N_31813 : std_logic ;
  signal N_31809 : std_logic ;
  signal N_31808 : std_logic ;
  signal N_31803 : std_logic ;
  signal N_31769 : std_logic ;
  signal N_31768 : std_logic ;
  signal N_31767 : std_logic ;
  signal N_31743 : std_logic ;
  signal N_31719 : std_logic ;
  signal N_31716 : std_logic ;
  signal N_31703 : std_logic ;
  signal N_31704 : std_logic ;
  signal N_31709 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1786\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2652\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1810\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2494\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2490\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2508\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2513\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8994\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_334\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2485\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1922\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1932\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1957\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2636\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2042\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2484\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2063\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2114\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2654\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2273\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2499\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2546\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2283\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2291\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2292\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2658\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2300\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2505\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_885_I\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2525\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2536\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2703\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2538\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2648\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2355\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2598\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_729\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_647\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2369\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2370\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2419\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2526\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2420\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2421\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2462\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2474\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2544\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2579\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2590\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2551\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2609\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2640\ : std_logic ;
  signal \GRLFPC2_0.N_38\ : std_logic ;
  signal \GRLFPC2_0.N_909_7\ : std_logic ;
  signal \GRLFPC2_0.N_94\ : std_logic ;
  signal \GRLFPC2_0.N_40\ : std_logic ;
  signal \GRLFPC2_0.N_78\ : std_logic ;
  signal \GRLFPC2_0.N_908_7\ : std_logic ;
  signal \GRLFPC2_0.N_77\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1902\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2337\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2341\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1816\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1819\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1815\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1811\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1812\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_568\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1808\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_450\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1042\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8639\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1940\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2263\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2127\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2639\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2342\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_726\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_354\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2214\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1969\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2422\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2572\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_318\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1164\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3942\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1903\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2354\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2351\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1982\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8695\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2290\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2288\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2274\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2268\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2267\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2581\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2534\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2373\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9074\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9074_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2302\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_445\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2586\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8752\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2587\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9079\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2367\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2784\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1954\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1967\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2311\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2306\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2405\ : std_logic ;
  signal N_33055 : std_logic ;
  signal N_33043_I : std_logic ;
  signal N_31887 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2504\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2762\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1967_1\ : std_logic ;
  signal N_28952 : std_logic ;
  signal N_28951 : std_logic ;
  signal N_28947 : std_logic ;
  signal N_28945 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2655\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2634\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2776\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2763\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2602\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2725\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2671\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2779\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_346\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2518\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_339\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2457\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2697\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2788\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2767\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2722\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2707\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2693\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2689\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2666\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2663\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2657\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2633\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MAPMULXFF.UN7_UNIMPMAP\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5771\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_12239\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_2_1_CO1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_12247\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1281_I\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10635\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6961\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_60.Z_1_CO0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_60.Z_1_CO1\ : std_logic ;
  signal N_34177 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3848\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7144\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4534\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3639\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\ : std_logic ;
  signal N_29788 : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_1\ : std_logic ;
  signal \GRLFPC2_0.N_1072_M\ : std_logic ;
  signal \GRLFPC2_0.COMB.RS1V_1\ : std_logic ;
  signal \GRLFPC2_0.N_2989\ : std_logic ;
  signal \GRLFPC2_0.N_2992\ : std_logic ;
  signal \GRLFPC2_0.N_2990\ : std_logic ;
  signal \GRLFPC2_0.N_2993\ : std_logic ;
  signal N_36304 : std_logic ;
  signal \GRLFPC2_0.N_2991\ : std_logic ;
  signal \GRLFPC2_0.RS1D_CNST\ : std_logic ;
  signal \GRLFPC2_0.COMB.FPDECODE.RDD6\ : std_logic ;
  signal \GRLFPC2_0.RS1V_0_SQMUXA_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.GEN\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5322\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5452\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7210\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5446\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN7_STKGEN\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_1_CO0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_947_I\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_959_I\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5324\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN25_GEN\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN13_GEN\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6583\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7782_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10013\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4662\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4233\ : std_logic ;
  signal \GRLFPC2_0.FPO.SIGN\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN1_R.I.V_1\ : std_logic ;
  signal \GRLFPC2_0.N_3422\ : std_logic ;
  signal \GRLFPC2_0.COMB.ISFPOP2_1\ : std_logic ;
  signal \GRLFPC2_0.COMB.ANNULRES_1\ : std_logic ;
  signal \GRLFPC2_0.N_1768\ : std_logic ;
  signal \GRLFPC2_0.N_158\ : std_logic ;
  signal \GRLFPC2_0.R.MK.RST_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TEMP\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10866\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10867\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10939\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10880\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10936\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10937\ : std_logic ;
  signal \GRLFPC2_0.N_3168\ : std_logic ;
  signal \GRLFPC2_0.N_1721\ : std_logic ;
  signal \GRLFPC2_0.N_1309\ : std_logic ;
  signal \GRLFPC2_0.V.FSR.CEXC_3_SQMUXA_1\ : std_logic ;
  signal \GRLFPC2_0.N_1586\ : std_logic ;
  signal \GRLFPC2_0.N_1515\ : std_logic ;
  signal \GRLFPC2_0.N_1302\ : std_logic ;
  signal \GRLFPC2_0.WREN2_2_SQMUXA\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_237\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10526\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10532\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10535\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10536\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10513\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10517\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10529\ : std_logic ;
  signal \GRLFPC2_0.N_3033\ : std_logic ;
  signal \GRLFPC2_0.N_3027\ : std_logic ;
  signal \GRLFPC2_0.N_3220\ : std_logic ;
  signal \GRLFPC2_0.N_3219\ : std_logic ;
  signal \GRLFPC2_0.N_3141\ : std_logic ;
  signal \GRLFPC2_0.R.I.V_1_0_G2\ : std_logic ;
  signal \GRLFPC2_0.N_3163\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10533\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10530\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10525\ : std_logic ;
  signal \GRLFPC2_0.N_3140\ : std_logic ;
  signal \GRLFPC2_0.N_145\ : std_logic ;
  signal \GRLFPC2_0.N_146\ : std_logic ;
  signal \GRLFPC2_0.N_3144\ : std_logic ;
  signal \GRLFPC2_0.N_3145\ : std_logic ;
  signal \GRLFPC2_0.N_3146\ : std_logic ;
  signal \GRLFPC2_0.N_3147\ : std_logic ;
  signal \GRLFPC2_0.N_151\ : std_logic ;
  signal \GRLFPC2_0.N_152\ : std_logic ;
  signal \GRLFPC2_0.N_153\ : std_logic ;
  signal \GRLFPC2_0.N_3151\ : std_logic ;
  signal \GRLFPC2_0.N_3152\ : std_logic ;
  signal \GRLFPC2_0.N_156\ : std_logic ;
  signal \GRLFPC2_0.N_157\ : std_logic ;
  signal \GRLFPC2_0.N_3122\ : std_logic ;
  signal \GRLFPC2_0.N_3156\ : std_logic ;
  signal \GRLFPC2_0.N_3125\ : std_logic ;
  signal \GRLFPC2_0.N_3160\ : std_logic ;
  signal \GRLFPC2_0.N_3128\ : std_logic ;
  signal \GRLFPC2_0.N_3162\ : std_logic ;
  signal \GRLFPC2_0.N_3164\ : std_logic ;
  signal \GRLFPC2_0.N_3165\ : std_logic ;
  signal \GRLFPC2_0.N_3134\ : std_logic ;
  signal \GRLFPC2_0.N_3136\ : std_logic ;
  signal \GRLFPC2_0.N_141\ : std_logic ;
  signal \GRLFPC2_0.N_140\ : std_logic ;
  signal \GRLFPC2_0.N_3429\ : std_logic ;
  signal \GRLFPC2_0.N_3428\ : std_logic ;
  signal \GRLFPC2_0.N_3427\ : std_logic ;
  signal \GRLFPC2_0.N_3426\ : std_logic ;
  signal \GRLFPC2_0.N_3227\ : std_logic ;
  signal \GRLFPC2_0.N_3226\ : std_logic ;
  signal \GRLFPC2_0.N_3032\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9989\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10016\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9829\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9978\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10211\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9797\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.UN17_U_RDN\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10007\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10006\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10010\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10015\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10870\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10883\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10003\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9790\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9833\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9975\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9993\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10210\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10209\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10208\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9994\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9983\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9972\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9971\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9970\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9997\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9968\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9996\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9979\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9995\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9998\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9844\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10000\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9999\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9789\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9981\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9985\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10008\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10011\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10884\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10017\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10018\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10206\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9992\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9986\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10019\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9984\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10207\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10205\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9969\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9791\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9990\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9982\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9980\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9828\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10001\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10002\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9974\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9991\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9987\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9988\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9976\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9977\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10012\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10014\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10634\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10944\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10935\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10872\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10886\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10869\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10882\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10868\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10881\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10879\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10865\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10878\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10890\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10887\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10885\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10889\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10888\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10520\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10514\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10579\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10553\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10554\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN11_WQSTSETS\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7035\ : std_logic ;
  signal \GRLFPC2_0.N_10\ : std_logic ;
  signal \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA\ : std_logic ;
  signal \GRLFPC2_0.N_11\ : std_logic ;
  signal \GRLFPC2_0.N_7\ : std_logic ;
  signal \GRLFPC2_0.N_1675_1\ : std_logic ;
  signal \GRLFPC2_0.N_1213\ : std_logic ;
  signal \GRLFPC2_0.N_1720\ : std_logic ;
  signal \GRLFPC2_0.N_2888\ : std_logic ;
  signal \GRLFPC2_0.N_1676\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1919\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_529\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN17_SHDVAR\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4664\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN18_XZXBUS_14\ : std_logic ;
  signal \GRLFPC2_0.N_1669\ : std_logic ;
  signal \GRLFPC2_0.V.FSR.FTT_1_SQMUXA_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2726\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_329\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2757\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7051\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7034\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5339\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5343\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5301\ : std_logic ;
  signal N_52211 : std_logic ;
  signal N_52474 : std_logic ;
  signal N_52547 : std_logic ;
  signal N_52556 : std_logic ;
  signal N_52645 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_A3_0_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O2_1\ : std_logic ;
  signal N_52547_TZ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_3\ : std_logic ;
  signal N_55054 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN10_FEEDBACK\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_12_TZ\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_1_TZ\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_13_TZ\ : std_logic ;
  signal \GRLFPC2_0.WREN2_1_SQMUXA_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_27_S_0\ : std_logic ;
  signal N_32052_1 : std_logic ;
  signal N_33133_1 : std_logic ;
  signal N_33069 : std_logic ;
  signal N_32159 : std_logic ;
  signal N_31921_3 : std_logic ;
  signal N_31924_1 : std_logic ;
  signal N_31925_1 : std_logic ;
  signal \GRLFPC2_0.N_27\ : std_logic ;
  signal N_32243 : std_logic ;
  signal \GRLFPC2_0.R.A.LD_0_0_G1_0\ : std_logic ;
  signal \GRLFPC2_0.V.FSR.CEXC_2_SQMUXA_0\ : std_logic ;
  signal N_57352 : std_logic ;
  signal N_57353 : std_logic ;
  signal N_57354 : std_logic ;
  signal N_57355 : std_logic ;
  signal N_57356 : std_logic ;
  signal N_57357 : std_logic ;
  signal N_57358 : std_logic ;
  signal N_57359 : std_logic ;
  signal N_57360 : std_logic ;
  signal N_57361 : std_logic ;
  signal N_57362 : std_logic ;
  signal N_57363 : std_logic ;
  signal N_57364 : std_logic ;
  signal N_57365 : std_logic ;
  signal N_57366 : std_logic ;
  signal N_57367 : std_logic ;
  signal N_57368 : std_logic ;
  signal N_57369 : std_logic ;
  signal N_57370 : std_logic ;
  signal N_57371 : std_logic ;
  signal N_57372 : std_logic ;
  signal N_57373 : std_logic ;
  signal N_57374 : std_logic ;
  signal N_57375 : std_logic ;
  signal N_57376 : std_logic ;
  signal N_57377 : std_logic ;
  signal N_57378 : std_logic ;
  signal N_57379 : std_logic ;
  signal N_57380 : std_logic ;
  signal N_57381 : std_logic ;
  signal N_57382 : std_logic ;
  signal N_57383 : std_logic ;
  signal N_57384 : std_logic ;
  signal N_57385 : std_logic ;
  signal N_57386 : std_logic ;
  signal N_57387 : std_logic ;
  signal N_57388 : std_logic ;
  signal N_57389 : std_logic ;
  signal N_57392 : std_logic ;
  signal N_57393 : std_logic ;
  signal N_57394 : std_logic ;
  signal N_57395 : std_logic ;
  signal N_57396 : std_logic ;
  signal N_57397 : std_logic ;
  signal N_57398 : std_logic ;
  signal N_57399 : std_logic ;
  signal N_57400 : std_logic ;
  signal N_57401 : std_logic ;
  signal N_57402 : std_logic ;
  signal N_57403 : std_logic ;
  signal N_57404 : std_logic ;
  signal N_57405 : std_logic ;
  signal N_57406 : std_logic ;
  signal N_57407 : std_logic ;
  signal N_57408 : std_logic ;
  signal N_57409 : std_logic ;
  signal N_57410 : std_logic ;
  signal N_57411 : std_logic ;
  signal N_57412 : std_logic ;
  signal N_57413 : std_logic ;
  signal N_57414 : std_logic ;
  signal N_57415 : std_logic ;
  signal N_57416 : std_logic ;
  signal N_57417 : std_logic ;
  signal N_57418 : std_logic ;
  signal N_57419 : std_logic ;
  signal N_57420 : std_logic ;
  signal N_57421 : std_logic ;
  signal N_57422 : std_logic ;
  signal N_57423 : std_logic ;
  signal N_57424 : std_logic ;
  signal N_57425 : std_logic ;
  signal N_57426 : std_logic ;
  signal N_57427 : std_logic ;
  signal N_57428 : std_logic ;
  signal N_57429 : std_logic ;
  signal N_57430 : std_logic ;
  signal N_57431 : std_logic ;
  signal N_57432 : std_logic ;
  signal N_57433 : std_logic ;
  signal N_57434 : std_logic ;
  signal N_57435 : std_logic ;
  signal N_57436 : std_logic ;
  signal N_57437 : std_logic ;
  signal N_57438 : std_logic ;
  signal N_57439 : std_logic ;
  signal N_57440 : std_logic ;
  signal N_57441 : std_logic ;
  signal N_57442 : std_logic ;
  signal N_57443 : std_logic ;
  signal N_57444 : std_logic ;
  signal N_57445 : std_logic ;
  signal N_57446 : std_logic ;
  signal N_57447 : std_logic ;
  signal N_57448 : std_logic ;
  signal N_57449 : std_logic ;
  signal N_57450 : std_logic ;
  signal N_57451 : std_logic ;
  signal N_57452 : std_logic ;
  signal N_57453 : std_logic ;
  signal N_57454 : std_logic ;
  signal N_57455 : std_logic ;
  signal N_57456 : std_logic ;
  signal N_57457 : std_logic ;
  signal N_57458 : std_logic ;
  signal N_57459 : std_logic ;
  signal N_57460 : std_logic ;
  signal N_57461 : std_logic ;
  signal N_57462 : std_logic ;
  signal N_57463 : std_logic ;
  signal N_57464 : std_logic ;
  signal N_57465 : std_logic ;
  signal N_57466 : std_logic ;
  signal N_57467 : std_logic ;
  signal N_57468 : std_logic ;
  signal N_57469 : std_logic ;
  signal N_57470 : std_logic ;
  signal N_57471 : std_logic ;
  signal N_57472 : std_logic ;
  signal N_57473 : std_logic ;
  signal N_57474 : std_logic ;
  signal N_57475 : std_logic ;
  signal N_57476 : std_logic ;
  signal N_57477 : std_logic ;
  signal N_57478 : std_logic ;
  signal N_57479 : std_logic ;
  signal N_57480 : std_logic ;
  signal N_57481 : std_logic ;
  signal N_57482 : std_logic ;
  signal N_57483 : std_logic ;
  signal N_57484 : std_logic ;
  signal N_57485 : std_logic ;
  signal N_57486 : std_logic ;
  signal N_57487 : std_logic ;
  signal N_57488 : std_logic ;
  signal N_57489 : std_logic ;
  signal N_57490 : std_logic ;
  signal N_57491 : std_logic ;
  signal N_57492 : std_logic ;
  signal N_57493 : std_logic ;
  signal N_57494 : std_logic ;
  signal N_57495 : std_logic ;
  signal N_57496 : std_logic ;
  signal N_57497 : std_logic ;
  signal N_57498 : std_logic ;
  signal N_57499 : std_logic ;
  signal N_57500 : std_logic ;
  signal N_57501 : std_logic ;
  signal N_57502 : std_logic ;
  signal N_57503 : std_logic ;
  signal N_57504 : std_logic ;
  signal N_57505 : std_logic ;
  signal N_57506 : std_logic ;
  signal N_57507 : std_logic ;
  signal N_57508 : std_logic ;
  signal N_57509 : std_logic ;
  signal N_57510 : std_logic ;
  signal N_57511 : std_logic ;
  signal N_57512 : std_logic ;
  signal N_57513 : std_logic ;
  signal N_57514 : std_logic ;
  signal N_57515 : std_logic ;
  signal N_57516 : std_logic ;
  signal N_57517 : std_logic ;
  signal N_57518 : std_logic ;
  signal N_57519 : std_logic ;
  signal N_57520 : std_logic ;
  signal N_57521 : std_logic ;
  signal N_57522 : std_logic ;
  signal N_57523 : std_logic ;
  signal N_57524 : std_logic ;
  signal N_57525 : std_logic ;
  signal N_57526 : std_logic ;
  signal N_57527 : std_logic ;
  signal N_57528 : std_logic ;
  signal N_57529 : std_logic ;
  signal N_57530 : std_logic ;
  signal N_57531 : std_logic ;
  signal N_57532 : std_logic ;
  signal N_57533 : std_logic ;
  signal N_57534 : std_logic ;
  signal N_57535 : std_logic ;
  signal N_57536 : std_logic ;
  signal N_57537 : std_logic ;
  signal N_57538 : std_logic ;
  signal N_57539 : std_logic ;
  signal N_57540 : std_logic ;
  signal N_57541 : std_logic ;
  signal N_57542 : std_logic ;
  signal N_57543 : std_logic ;
  signal N_57544 : std_logic ;
  signal N_57545 : std_logic ;
  signal N_57546 : std_logic ;
  signal N_57547 : std_logic ;
  signal N_57548 : std_logic ;
  signal N_57549 : std_logic ;
  signal N_57550 : std_logic ;
  signal N_57551 : std_logic ;
  signal N_57552 : std_logic ;
  signal N_57553 : std_logic ;
  signal N_57554 : std_logic ;
  signal N_57555 : std_logic ;
  signal N_57556 : std_logic ;
  signal N_57557 : std_logic ;
  signal N_57558 : std_logic ;
  signal N_57559 : std_logic ;
  signal N_57560 : std_logic ;
  signal N_57561 : std_logic ;
  signal N_57562 : std_logic ;
  signal N_57563 : std_logic ;
  signal N_57564 : std_logic ;
  signal N_57565 : std_logic ;
  signal N_57566 : std_logic ;
  signal N_57567 : std_logic ;
  signal N_57571 : std_logic ;
  signal N_57572 : std_logic ;
  signal N_57578 : std_logic ;
  signal N_57579 : std_logic ;
  signal N_57587 : std_logic ;
  signal N_57594 : std_logic ;
  signal N_57595 : std_logic ;
  signal N_57601 : std_logic ;
  signal N_57602 : std_logic ;
  signal N_57610 : std_logic ;
  signal N_57617 : std_logic ;
  signal N_57618 : std_logic ;
  signal N_57624 : std_logic ;
  signal N_57625 : std_logic ;
  signal N_57633 : std_logic ;
  signal N_57640 : std_logic ;
  signal N_57641 : std_logic ;
  signal N_57647 : std_logic ;
  signal N_57648 : std_logic ;
  signal N_57656 : std_logic ;
  signal N_57663 : std_logic ;
  signal N_57664 : std_logic ;
  signal N_57670 : std_logic ;
  signal N_57671 : std_logic ;
  signal N_57679 : std_logic ;
  signal N_57686 : std_logic ;
  signal N_57687 : std_logic ;
  signal N_57693 : std_logic ;
  signal N_57694 : std_logic ;
  signal N_57702 : std_logic ;
  signal N_57709 : std_logic ;
  signal N_57710 : std_logic ;
  signal N_57716 : std_logic ;
  signal N_57717 : std_logic ;
  signal N_57725 : std_logic ;
  signal N_57732 : std_logic ;
  signal N_57733 : std_logic ;
  signal N_57739 : std_logic ;
  signal N_57740 : std_logic ;
  signal N_57748 : std_logic ;
  signal N_57755 : std_logic ;
  signal N_57756 : std_logic ;
  signal N_57762 : std_logic ;
  signal N_57763 : std_logic ;
  signal N_57771 : std_logic ;
  signal N_57778 : std_logic ;
  signal N_57779 : std_logic ;
  signal N_57785 : std_logic ;
  signal N_57786 : std_logic ;
  signal N_57794 : std_logic ;
  signal N_57801 : std_logic ;
  signal N_57802 : std_logic ;
  signal N_57808 : std_logic ;
  signal N_57809 : std_logic ;
  signal N_57817 : std_logic ;
  signal N_57824 : std_logic ;
  signal N_57825 : std_logic ;
  signal N_57831 : std_logic ;
  signal N_57832 : std_logic ;
  signal N_57840 : std_logic ;
  signal N_57847 : std_logic ;
  signal N_57848 : std_logic ;
  signal N_57854 : std_logic ;
  signal N_57855 : std_logic ;
  signal N_57863 : std_logic ;
  signal N_57870 : std_logic ;
  signal N_57871 : std_logic ;
  signal N_57877 : std_logic ;
  signal N_57878 : std_logic ;
  signal N_57886 : std_logic ;
  signal N_57893 : std_logic ;
  signal N_57894 : std_logic ;
  signal N_57900 : std_logic ;
  signal N_57901 : std_logic ;
  signal N_57909 : std_logic ;
  signal N_57916 : std_logic ;
  signal N_57917 : std_logic ;
  signal N_57923 : std_logic ;
  signal N_57924 : std_logic ;
  signal N_57932 : std_logic ;
  signal N_57939 : std_logic ;
  signal N_57940 : std_logic ;
  signal N_57946 : std_logic ;
  signal N_57947 : std_logic ;
  signal N_57955 : std_logic ;
  signal N_57962 : std_logic ;
  signal N_57963 : std_logic ;
  signal N_57969 : std_logic ;
  signal N_57970 : std_logic ;
  signal N_57978 : std_logic ;
  signal N_57985 : std_logic ;
  signal N_57986 : std_logic ;
  signal N_57992 : std_logic ;
  signal N_57993 : std_logic ;
  signal N_58001 : std_logic ;
  signal N_58008 : std_logic ;
  signal N_58009 : std_logic ;
  signal N_58015 : std_logic ;
  signal N_58016 : std_logic ;
  signal N_58024 : std_logic ;
  signal N_58031 : std_logic ;
  signal N_58032 : std_logic ;
  signal N_58038 : std_logic ;
  signal N_58039 : std_logic ;
  signal N_58047 : std_logic ;
  signal N_58054 : std_logic ;
  signal N_58055 : std_logic ;
  signal N_58061 : std_logic ;
  signal N_58062 : std_logic ;
  signal N_58070 : std_logic ;
  signal N_58077 : std_logic ;
  signal N_58078 : std_logic ;
  signal N_58084 : std_logic ;
  signal N_58085 : std_logic ;
  signal N_58093 : std_logic ;
  signal N_58100 : std_logic ;
  signal N_58101 : std_logic ;
  signal N_58107 : std_logic ;
  signal N_58108 : std_logic ;
  signal N_58116 : std_logic ;
  signal N_58123 : std_logic ;
  signal N_58124 : std_logic ;
  signal N_58130 : std_logic ;
  signal N_58131 : std_logic ;
  signal N_58139 : std_logic ;
  signal N_58146 : std_logic ;
  signal N_58147 : std_logic ;
  signal N_58153 : std_logic ;
  signal N_58154 : std_logic ;
  signal N_58162 : std_logic ;
  signal N_58169 : std_logic ;
  signal N_58170 : std_logic ;
  signal N_58176 : std_logic ;
  signal N_58177 : std_logic ;
  signal N_58185 : std_logic ;
  signal N_58192 : std_logic ;
  signal N_58193 : std_logic ;
  signal N_58199 : std_logic ;
  signal N_58200 : std_logic ;
  signal N_58208 : std_logic ;
  signal N_58215 : std_logic ;
  signal N_58216 : std_logic ;
  signal N_58222 : std_logic ;
  signal N_58223 : std_logic ;
  signal N_58231 : std_logic ;
  signal N_58238 : std_logic ;
  signal N_58239 : std_logic ;
  signal N_58245 : std_logic ;
  signal N_58246 : std_logic ;
  signal N_58254 : std_logic ;
  signal N_58261 : std_logic ;
  signal N_58262 : std_logic ;
  signal N_58268 : std_logic ;
  signal N_58269 : std_logic ;
  signal N_58277 : std_logic ;
  signal N_58284 : std_logic ;
  signal N_58285 : std_logic ;
  signal N_58291 : std_logic ;
  signal N_58292 : std_logic ;
  signal N_58300 : std_logic ;
  signal N_58307 : std_logic ;
  signal N_58308 : std_logic ;
  signal N_58314 : std_logic ;
  signal N_58315 : std_logic ;
  signal N_58323 : std_logic ;
  signal N_58330 : std_logic ;
  signal N_58331 : std_logic ;
  signal N_58337 : std_logic ;
  signal N_58338 : std_logic ;
  signal N_58346 : std_logic ;
  signal N_58353 : std_logic ;
  signal N_58354 : std_logic ;
  signal N_58360 : std_logic ;
  signal N_58361 : std_logic ;
  signal N_58369 : std_logic ;
  signal N_58376 : std_logic ;
  signal N_58377 : std_logic ;
  signal N_58383 : std_logic ;
  signal N_58384 : std_logic ;
  signal N_58392 : std_logic ;
  signal N_58399 : std_logic ;
  signal N_58400 : std_logic ;
  signal N_58406 : std_logic ;
  signal N_58407 : std_logic ;
  signal N_58415 : std_logic ;
  signal N_58422 : std_logic ;
  signal N_58423 : std_logic ;
  signal N_58429 : std_logic ;
  signal N_58430 : std_logic ;
  signal N_58438 : std_logic ;
  signal N_58445 : std_logic ;
  signal N_58446 : std_logic ;
  signal N_58452 : std_logic ;
  signal N_58453 : std_logic ;
  signal N_58461 : std_logic ;
  signal N_58468 : std_logic ;
  signal N_58469 : std_logic ;
  signal N_58475 : std_logic ;
  signal N_58476 : std_logic ;
  signal N_58484 : std_logic ;
  signal N_58491 : std_logic ;
  signal N_58492 : std_logic ;
  signal N_58498 : std_logic ;
  signal N_58499 : std_logic ;
  signal N_58507 : std_logic ;
  signal N_58514 : std_logic ;
  signal N_58515 : std_logic ;
  signal N_58521 : std_logic ;
  signal N_58522 : std_logic ;
  signal N_58530 : std_logic ;
  signal N_58537 : std_logic ;
  signal N_58538 : std_logic ;
  signal N_58544 : std_logic ;
  signal N_58545 : std_logic ;
  signal N_58553 : std_logic ;
  signal N_58560 : std_logic ;
  signal N_58561 : std_logic ;
  signal N_58567 : std_logic ;
  signal N_58568 : std_logic ;
  signal N_58576 : std_logic ;
  signal N_58585 : std_logic ;
  signal N_58586 : std_logic ;
  signal N_58592 : std_logic ;
  signal N_58593 : std_logic ;
  signal N_58601 : std_logic ;
  signal N_58608 : std_logic ;
  signal N_58609 : std_logic ;
  signal N_58615 : std_logic ;
  signal N_58616 : std_logic ;
  signal N_58624 : std_logic ;
  signal N_58631 : std_logic ;
  signal N_58632 : std_logic ;
  signal N_58638 : std_logic ;
  signal N_58639 : std_logic ;
  signal N_58647 : std_logic ;
  signal N_58657 : std_logic ;
  signal N_58667 : std_logic ;
  signal N_58668 : std_logic ;
  signal N_58671 : std_logic ;
  signal N_58672 : std_logic ;
  signal N_58676 : std_logic ;
  signal N_58677 : std_logic ;
  signal N_58683 : std_logic ;
  signal N_58684 : std_logic ;
  signal N_58692 : std_logic ;
  signal N_58699 : std_logic ;
  signal N_58700 : std_logic ;
  signal N_58706 : std_logic ;
  signal N_58707 : std_logic ;
  signal N_58715 : std_logic ;
  signal N_58722 : std_logic ;
  signal N_58723 : std_logic ;
  signal N_58729 : std_logic ;
  signal N_58730 : std_logic ;
  signal N_58738 : std_logic ;
  signal N_58745 : std_logic ;
  signal N_58746 : std_logic ;
  signal N_58752 : std_logic ;
  signal N_58753 : std_logic ;
  signal N_58761 : std_logic ;
  signal N_58820 : std_logic ;
  signal N_58821 : std_logic ;
  signal N_58827 : std_logic ;
  signal N_58828 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3729_I_0\ : std_logic ;
  signal CPI_D_INST_INTERNAL_6 : std_logic ;
  signal \GRLFPC2_0.N_1830_O\ : std_logic ;
  signal \GRLFPC2_0.N_1683\ : std_logic ;
  signal \GRLFPC2_0.N_1237\ : std_logic ;
  signal \GRLFPC2_0.COMB.LOCKGEN.LOCKI_I_1\ : std_logic ;
  signal N_59162 : std_logic ;
  signal N_59163 : std_logic ;
  signal N_59164 : std_logic ;
  signal N_59166 : std_logic ;
  signal N_59168 : std_logic ;
  signal N_59169 : std_logic ;
  signal N_59170 : std_logic ;
  signal N_59171 : std_logic ;
  signal N_59172 : std_logic ;
  signal N_59173 : std_logic ;
  signal N_59174 : std_logic ;
  signal N_59178 : std_logic ;
  signal N_59179 : std_logic ;
  signal N_59180 : std_logic ;
  signal N_59183 : std_logic ;
  signal N_59185 : std_logic ;
  signal N_59186 : std_logic ;
  signal N_59187 : std_logic ;
  signal N_59188 : std_logic ;
  signal N_59189 : std_logic ;
  signal N_59191 : std_logic ;
  signal N_59192 : std_logic ;
  signal N_59193 : std_logic ;
  signal N_59194 : std_logic ;
  signal N_59195 : std_logic ;
  signal N_59196 : std_logic ;
  signal N_59197 : std_logic ;
  signal N_59199 : std_logic ;
  signal N_59200 : std_logic ;
  signal N_59205 : std_logic ;
  signal N_59206 : std_logic ;
  signal N_59208 : std_logic ;
  signal N_59209 : std_logic ;
  signal N_59210 : std_logic ;
  signal N_59211 : std_logic ;
  signal N_59213 : std_logic ;
  signal N_59215 : std_logic ;
  signal N_59217 : std_logic ;
  signal N_59218 : std_logic ;
  signal N_59219 : std_logic ;
  signal N_59220 : std_logic ;
  signal N_59226 : std_logic ;
  signal N_59228 : std_logic ;
  signal N_59229 : std_logic ;
  signal N_59232 : std_logic ;
  signal N_59234 : std_logic ;
  signal N_59235 : std_logic ;
  signal N_59236 : std_logic ;
  signal N_59237 : std_logic ;
  signal N_59238 : std_logic ;
  signal N_59239 : std_logic ;
  signal N_59240 : std_logic ;
  signal N_59242 : std_logic ;
  signal N_59243 : std_logic ;
  signal N_59244 : std_logic ;
  signal N_59245 : std_logic ;
  signal N_59246 : std_logic ;
  signal N_59249 : std_logic ;
  signal N_59250 : std_logic ;
  signal N_59251 : std_logic ;
  signal N_59252 : std_logic ;
  signal N_59253 : std_logic ;
  signal N_59254 : std_logic ;
  signal N_59255 : std_logic ;
  signal N_59258 : std_logic ;
  signal N_59260 : std_logic ;
  signal N_59261 : std_logic ;
  signal N_59262 : std_logic ;
  signal N_59263 : std_logic ;
  signal N_59264 : std_logic ;
  signal N_59265 : std_logic ;
  signal N_59267 : std_logic ;
  signal N_59268 : std_logic ;
  signal N_59269 : std_logic ;
  signal N_59270 : std_logic ;
  signal N_59271 : std_logic ;
  signal N_59272 : std_logic ;
  signal N_59273 : std_logic ;
  signal N_59274 : std_logic ;
  signal N_59275 : std_logic ;
  signal N_59281 : std_logic ;
  signal N_59283 : std_logic ;
  signal N_59284 : std_logic ;
  signal N_59285 : std_logic ;
  signal N_59286 : std_logic ;
  signal N_59287 : std_logic ;
  signal N_59288 : std_logic ;
  signal N_59291 : std_logic ;
  signal N_59293 : std_logic ;
  signal N_59294 : std_logic ;
  signal N_59297 : std_logic ;
  signal N_59304 : std_logic ;
  signal N_59307 : std_logic ;
  signal N_59308 : std_logic ;
  signal N_59309 : std_logic ;
  signal N_59311 : std_logic ;
  signal N_59317 : std_logic ;
  signal N_59318 : std_logic ;
  signal N_59319 : std_logic ;
  signal N_59323 : std_logic ;
  signal N_59328 : std_logic ;
  signal N_59331 : std_logic ;
  signal N_59336 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_15_TZ\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_1_TZ\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_6_TZ\ : std_logic ;
  signal \GRLFPC2_0.COMB.WREN2_9_IV_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.WREN2_9_IV_1\ : std_logic ;
  signal \GRLFPC2_0.COMB.WREN1_9_IV_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.WREN1_9_IV_1\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN8_CCV_2\ : std_logic ;
  signal \GRLFPC2_0.COMB.RDD_1.M14_0_A2_3\ : std_logic ;
  signal \GRLFPC2_0.COMB.FPDECODE.UN1_FPCI_7_4\ : std_logic ;
  signal \GRLFPC2_0.COMB.SEQERR.UN13_OP_0_3\ : std_logic ;
  signal \GRLFPC2_0.UN1_MOV_1_SQMUXA_0\ : std_logic ;
  signal \GRLFPC2_0.MOV_2_SQMUXA_1\ : std_logic ;
  signal \GRLFPC2_0.COMB.RSDECODE.UN1_FPCI_1\ : std_logic ;
  signal \GRLFPC2_0.COMB.RSDECODE.UN1_FPCI_2\ : std_logic ;
  signal \GRLFPC2_0.ANNULRES_0_SQMUXA_10_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.A.SEQERR_1_0_A2_0_3\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN1_MEXC_1_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN1_MEXC_1_1\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN1_FPCI_3_1\ : std_logic ;
  signal \GRLFPC2_0.COMB.ANNULFPU_1_U_0_0\ : std_logic ;
  signal \GRLFPC2_0.V.FSR.FTT_3_SQMUXA_I_A3_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4167_I_0_I_A3_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4167_I_0_I_A3_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN26_NOTAINFNAN_4\ : std_logic ;
  signal \GRLFPC2_0.COMB.ANNULRES_1_IV_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_4\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.A.RF2REN_1_0_7690_I_A5_0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7612_I_A7_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7612_I_A7_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7612_I_A7_10\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.A.RF1REN_1_0_7636_I_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_4914_1_A2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_19\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_20\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_22\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_23\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_26\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_27\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_28\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN2_HOLDN_0_A3_7\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN2_HOLDN_0_A3_8\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN2_HOLDN_0_A3_10\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN2_HOLDN_0_A3_11\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN2_HOLDN_0_A3_13\ : std_logic ;
  signal \GRLFPC2_0.R.E.AFSR_RET_0_0_G1_3\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN6_IUEXEC_1\ : std_logic ;
  signal \GRLFPC2_0.R.E.AFQ_RET_0_0_G1_4\ : std_logic ;
  signal \GRLFPC2_0.R.E.AFQ_RET_0_0_G1_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7612_I_1_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN12_SRTOSTICKY_3\ : std_logic ;
  signal \GRLFPC2_0.N_939_I_0_A2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_1__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_8__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_44__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_23__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_39__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_43__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_5_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_16\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_35__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_35__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_24__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_15_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_10_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_16\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_0_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_16\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_19\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_23\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_30__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_18\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_20\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_21\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1_0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_16__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_16__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_13_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_20\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_16\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_18\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_20\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_24\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_1_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.STARTSHFT.UN2_NOTDECODEDUNIMP_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_16\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_19\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_20\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_8\ : std_logic ;
  signal \GRLFPC2_0.R.I.V_1_0_G0_I_O4_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_16\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__G2_0_7242_I_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_242__G2_0_7304_I_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_243__G2_0_7273_I_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_241__G2_0_7335_I_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_19\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_21\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_23\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_25\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_27\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_31\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_32\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_36\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_37\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_38\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_39\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_40\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_42\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_45\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_46\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_49\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_50\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_52\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_53\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_240__G2_0_7366_I_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_239__G2_0_7397_I_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_238__G2_0_7428_I_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_237__G2_0_7459_I_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.MIFROMINST_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN30_CONDITIONAL_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.BUSYMULXFF.UN2_TEMP_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_I_0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2\ : std_logic ;
  signal \GRLFPC2_0.N_1470\ : std_logic ;
  signal \GRLFPC2_0.COMB.LOCKGEN.LOCKI_I_I\ : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\ : std_logic ;
  signal \GRLFPC2_0.WRADDR_0_SQMUXA_1\ : std_logic ;
  signal \GRLFPC2_0.N_1132\ : std_logic ;
  signal \GRLFPC2_0.V.FSR.CEXC_0_SQMUXA\ : std_logic ;
  signal \GRLFPC2_0.N_1517\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.E.STDATA2\ : std_logic ;
  signal \GRLFPC2_0.COMB.RDD_2\ : std_logic ;
  signal \GRLFPC2_0.N_1570\ : std_logic ;
  signal \GRLFPC2_0.N_1243\ : std_logic ;
  signal \GRLFPC2_0.WRADDR_1_SQMUXA\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.NOTPROP_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.NOTPROP\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10538\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2498\ : std_logic ;
  signal N_31921_1 : std_logic ;
  signal N_32141_1 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_255\ : std_logic ;
  signal N_31725_1 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\ : std_logic ;
  signal \GRLFPC2_0.N_1255\ : std_logic ;
  signal \GRLFPC2_0.R.I.EXC_2_0_4__N_5\ : std_logic ;
  signal N_76337 : std_logic ;
  signal \GRLFPC2_0.R.I.INST_1_0_9__G2\ : std_logic ;
  signal \GRLFPC2_0.R.A.AFSR\ : std_logic ;
  signal \GRLFPC2_0.R.A.AFQ\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422\ : std_logic ;
  signal N_76344 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN1_FPCI_4\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN1_R.A.RS1_1\ : std_logic ;
  signal N_79923 : std_logic ;
  signal N_79931 : std_logic ;
  signal N_79935 : std_logic ;
  signal N_79937 : std_logic ;
  signal N_79939 : std_logic ;
  signal N_79941 : std_logic ;
  signal N_79943 : std_logic ;
  signal N_79982 : std_logic ;
  signal N_79986 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5394\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349_I_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G0_0_O2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G1_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G0_I_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G0_I_0_2_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G0_I_0_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0_4__G0_4_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0_4__G0_2_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO\ : std_logic ;
  signal N_1_0 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2809_1_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_729_RETO\ : std_logic ;
  signal N_1_1 : std_logic ;
  signal N_28946_RETO : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_RETO\ : std_logic ;
  signal N_1_2 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO\ : std_logic ;
  signal N_1_3 : std_logic ;
  signal N_28947_RETO : std_logic ;
  signal N_1_4 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO\ : std_logic ;
  signal N_28945_RETO : std_logic ;
  signal N_1_5 : std_logic ;
  signal N_28950_RETO : std_logic ;
  signal N_1_6 : std_logic ;
  signal N_28951_RETO : std_logic ;
  signal N_1_7 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO\ : std_logic ;
  signal N_28952_RETO : std_logic ;
  signal N_1_8 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349_I_0_RETI\ : std_logic ;
  signal N_15 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5394_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2463_RETO\ : std_logic ;
  signal N_31763_1_RETO : std_logic ;
  signal N_31723_1_RETO : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_255_RETO\ : std_logic ;
  signal N_1_9 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_455_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2555_RETO\ : std_logic ;
  signal N_1_10 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_217_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2457_RETO\ : std_logic ;
  signal N_1_11 : std_logic ;
  signal RST_RETO : std_logic ;
  signal N_1_12 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO\ : std_logic ;
  signal N_1_13 : std_logic ;
  signal N_1_14 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I_RETO\ : std_logic ;
  signal N_1_15 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_RETO\ : std_logic ;
  signal N_1_16 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO\ : std_logic ;
  signal N_1_17 : std_logic ;
  signal N_80376 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.UN17_U_RDN_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.TEMP_RETO\ : std_logic ;
  signal N_1_18 : std_logic ;
  signal N_80377 : std_logic ;
  signal N_79941_RETO : std_logic ;
  signal N_1_19 : std_logic ;
  signal \GRLFPC2_0.FPO.BUSY_O\ : std_logic ;
  signal N_1_20 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3924_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.BUSYMULXFF.UN2_TEMP_2_RETO\ : std_logic ;
  signal N_1_21 : std_logic ;
  signal N_1_22 : std_logic ;
  signal N_1_23 : std_logic ;
  signal N_1_24 : std_logic ;
  signal N_1_25 : std_logic ;
  signal N_1_26 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO\ : std_logic ;
  signal N_1_27 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_319__G1_RETO\ : std_logic ;
  signal N_1_28 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_318__G1_RETO\ : std_logic ;
  signal N_1_29 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_372__G1_RETO\ : std_logic ;
  signal N_1_30 : std_logic ;
  signal N_1_31 : std_logic ;
  signal N_1_32 : std_logic ;
  signal N_1_33 : std_logic ;
  signal N_1_34 : std_logic ;
  signal N_1_35 : std_logic ;
  signal N_1_36 : std_logic ;
  signal N_1_37 : std_logic ;
  signal N_1_38 : std_logic ;
  signal N_1_39 : std_logic ;
  signal N_1_40 : std_logic ;
  signal N_1_41 : std_logic ;
  signal N_1_42 : std_logic ;
  signal N_1_43 : std_logic ;
  signal N_1_44 : std_logic ;
  signal N_1_45 : std_logic ;
  signal N_1_46 : std_logic ;
  signal N_1_47 : std_logic ;
  signal N_1_48 : std_logic ;
  signal N_1_49 : std_logic ;
  signal N_1_50 : std_logic ;
  signal N_1_51 : std_logic ;
  signal N_1_52 : std_logic ;
  signal N_1_53 : std_logic ;
  signal N_1_54 : std_logic ;
  signal N_1_55 : std_logic ;
  signal N_1_56 : std_logic ;
  signal N_1_57 : std_logic ;
  signal N_1_58 : std_logic ;
  signal N_1_59 : std_logic ;
  signal N_1_60 : std_logic ;
  signal N_1_61 : std_logic ;
  signal N_1_62 : std_logic ;
  signal N_1_63 : std_logic ;
  signal N_1_64 : std_logic ;
  signal N_1_65 : std_logic ;
  signal N_1_66 : std_logic ;
  signal N_1_67 : std_logic ;
  signal N_1_68 : std_logic ;
  signal N_1_69 : std_logic ;
  signal N_1_70 : std_logic ;
  signal N_1_71 : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_RETO\ : std_logic ;
  signal N_1_72 : std_logic ;
  signal N_1_73 : std_logic ;
  signal N_1_74 : std_logic ;
  signal N_1_75 : std_logic ;
  signal N_1_76 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO\ : std_logic ;
  signal N_1_77 : std_logic ;
  signal N_1_78 : std_logic ;
  signal N_1_79 : std_logic ;
  signal N_1_80 : std_logic ;
  signal N_1_81 : std_logic ;
  signal N_1_82 : std_logic ;
  signal N_1_83 : std_logic ;
  signal N_79998_RETO : std_logic ;
  signal N_1_84 : std_logic ;
  signal N_1_85 : std_logic ;
  signal N_1_86 : std_logic ;
  signal N_1_87 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G1_1_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_237_RETO\ : std_logic ;
  signal N_1_88 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2474_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1164_RETO\ : std_logic ;
  signal N_1_89 : std_logic ;
  signal N_1_90 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5330_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_I_0_0_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO\ : std_logic ;
  signal N_1_91 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_377_RETO\ : std_logic ;
  signal N_1_92 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO\ : std_logic ;
  signal N_1_93 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\ : std_logic ;
  signal N_28949_RETO : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO\ : std_logic ;
  signal N_1_94 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2466_1_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO\ : std_logic ;
  signal N_1_95 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10927_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_27_S_0_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10918_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO\ : std_logic ;
  signal N_55054_RETO : std_logic ;
  signal N_1_96 : std_logic ;
  signal N_26534_RETO : std_logic ;
  signal N_26560_RETO : std_logic ;
  signal N_26559_RETO : std_logic ;
  signal N_1_97 : std_logic ;
  signal N_26564_RETO : std_logic ;
  signal N_26563_RETO : std_logic ;
  signal N_1_98 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_175__G2_RETO\ : std_logic ;
  signal N_1_99 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_176__G2_RETO\ : std_logic ;
  signal N_1_100 : std_logic ;
  signal N_1_101 : std_logic ;
  signal N_1_102 : std_logic ;
  signal N_1_103 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_RETO\ : std_logic ;
  signal N_1_104 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_RETO\ : std_logic ;
  signal N_1_105 : std_logic ;
  signal N_1_106 : std_logic ;
  signal N_1_107 : std_logic ;
  signal N_1_108 : std_logic ;
  signal N_1_109 : std_logic ;
  signal N_1_110 : std_logic ;
  signal N_1_111 : std_logic ;
  signal N_1_112 : std_logic ;
  signal N_1_113 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2462_RETO\ : std_logic ;
  signal N_1_114 : std_logic ;
  signal N_80614 : std_logic ;
  signal N_80615 : std_logic ;
  signal N_80616 : std_logic ;
  signal N_80617 : std_logic ;
  signal N_80618 : std_logic ;
  signal N_80619 : std_logic ;
  signal N_80620 : std_logic ;
  signal N_80621 : std_logic ;
  signal N_80622 : std_logic ;
  signal N_80623 : std_logic ;
  signal N_80624 : std_logic ;
  signal N_80625 : std_logic ;
  signal N_80626 : std_logic ;
  signal N_80627 : std_logic ;
  signal N_80628 : std_logic ;
  signal N_80629 : std_logic ;
  signal N_80630 : std_logic ;
  signal N_80631 : std_logic ;
  signal N_80632 : std_logic ;
  signal N_80633 : std_logic ;
  signal N_80634 : std_logic ;
  signal N_80635 : std_logic ;
  signal N_80636 : std_logic ;
  signal N_80637 : std_logic ;
  signal N_80638 : std_logic ;
  signal N_80639 : std_logic ;
  signal N_80640 : std_logic ;
  signal N_80641 : std_logic ;
  signal N_80642 : std_logic ;
  signal N_80643 : std_logic ;
  signal N_80644 : std_logic ;
  signal N_80645 : std_logic ;
  signal N_80646 : std_logic ;
  signal N_80647 : std_logic ;
  signal N_80648 : std_logic ;
  signal N_80649 : std_logic ;
  signal N_80650 : std_logic ;
  signal N_80651 : std_logic ;
  signal N_80652 : std_logic ;
  signal N_80653 : std_logic ;
  signal N_80654 : std_logic ;
  signal N_80655 : std_logic ;
  signal N_80656 : std_logic ;
  signal N_80657 : std_logic ;
  signal N_80658 : std_logic ;
  signal N_80659 : std_logic ;
  signal N_80660 : std_logic ;
  signal N_80661 : std_logic ;
  signal N_80662 : std_logic ;
  signal N_80663 : std_logic ;
  signal N_80664 : std_logic ;
  signal N_80665 : std_logic ;
  signal N_80666 : std_logic ;
  signal N_80667 : std_logic ;
  signal N_80668 : std_logic ;
  signal N_80669 : std_logic ;
  signal N_80670 : std_logic ;
  signal N_80671 : std_logic ;
  signal N_80672 : std_logic ;
  signal N_80673 : std_logic ;
  signal N_80674 : std_logic ;
  signal N_81152 : std_logic ;
  signal N_81171 : std_logic ;
  signal N_81177 : std_logic ;
  signal N_81224 : std_logic ;
  signal N_81248 : std_logic ;
  signal N_81250 : std_logic ;
  signal N_81259 : std_logic ;
  signal N_81263 : std_logic ;
  signal N_81293 : std_logic ;
  signal N_81301 : std_logic ;
  signal N_81507 : std_logic ;
  signal N_81559 : std_logic ;
  signal N_81561 : std_logic ;
  signal N_81563 : std_logic ;
  signal N_81599 : std_logic ;
  signal N_81609 : std_logic ;
  signal N_81611 : std_logic ;
  signal N_81615 : std_logic ;
  signal N_81619 : std_logic ;
  signal N_81621 : std_logic ;
  signal N_81626 : std_logic ;
  signal N_81630 : std_logic ;
  signal N_81634 : std_logic ;
  signal N_81640 : std_logic ;
  signal N_81674 : std_logic ;
  signal N_81684 : std_logic ;
  signal N_81690 : std_logic ;
  signal N_81707 : std_logic ;
  signal N_81709 : std_logic ;
  signal N_81711 : std_logic ;
  signal N_81973 : std_logic ;
  signal N_81974 : std_logic ;
  signal N_81985 : std_logic ;
  signal N_81986 : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_I\ : std_logic ;
  signal N_26534_I : std_logic ;
  signal RST_I : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_RETI_0\ : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\ : std_logic ;
  signal N_32048_1_0 : std_logic ;
  signal N_32340_1_0 : std_logic ;
  signal N_31725_1_0 : std_logic ;
  signal N_31921_1_0 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10936_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10939_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10936_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10939_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10944_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10944_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4534_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897_0\ : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4534_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897_1\ : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10937_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10937_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN12_SRTOSTICKY_3_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G0_I_0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349_I_0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_0\ : std_logic ;
  signal N_28946_RETO_0 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_1\ : std_logic ;
  signal N_28946_RETO_1 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_2\ : std_logic ;
  signal N_28946_RETO_2 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_3\ : std_logic ;
  signal N_28946_RETO_3 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_RETO_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_4\ : std_logic ;
  signal N_28946_RETO_4 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_RETO_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_5\ : std_logic ;
  signal N_28946_RETO_5 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_RETO_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_6\ : std_logic ;
  signal N_28946_RETO_6 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_RETO_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_7\ : std_logic ;
  signal N_28946_RETO_7 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_RETO_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_16\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_16\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_17\ : std_logic ;
  signal N_28947_RETO_0 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_18\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_18\ : std_logic ;
  signal N_28947_RETO_1 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_19\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_19\ : std_logic ;
  signal N_28947_RETO_2 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_20\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_20\ : std_logic ;
  signal N_28947_RETO_3 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_21\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_21\ : std_logic ;
  signal N_28947_RETO_4 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_22\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_22\ : std_logic ;
  signal N_28947_RETO_5 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_23\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_23\ : std_logic ;
  signal N_28947_RETO_6 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_24\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_24\ : std_logic ;
  signal N_28947_RETO_7 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_25\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_25\ : std_logic ;
  signal N_28947_RETO_8 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_26\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_26\ : std_logic ;
  signal N_28947_RETO_9 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_27\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_27\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO_0\ : std_logic ;
  signal N_28945_RETO_0 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_28\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_28\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO_1\ : std_logic ;
  signal N_28945_RETO_1 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_29\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_29\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO_2\ : std_logic ;
  signal N_28945_RETO_2 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_30\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_30\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO_3\ : std_logic ;
  signal N_28945_RETO_3 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_31\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_31\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO_4\ : std_logic ;
  signal N_28945_RETO_4 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_32\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_32\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO_5\ : std_logic ;
  signal N_28945_RETO_5 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_33\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_33\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO_6\ : std_logic ;
  signal N_28945_RETO_6 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_34\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_34\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO_7\ : std_logic ;
  signal N_28945_RETO_7 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_35\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_35\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO_8\ : std_logic ;
  signal N_28945_RETO_8 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_36\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_36\ : std_logic ;
  signal N_28950_RETO_0 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_37\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_37\ : std_logic ;
  signal N_28950_RETO_1 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_38\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_38\ : std_logic ;
  signal N_28950_RETO_2 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_39\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_39\ : std_logic ;
  signal N_28950_RETO_3 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_40\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_40\ : std_logic ;
  signal N_28950_RETO_4 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_41\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_41\ : std_logic ;
  signal N_28950_RETO_5 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_42\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_42\ : std_logic ;
  signal N_28950_RETO_6 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_43\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_43\ : std_logic ;
  signal N_28950_RETO_7 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_44\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_44\ : std_logic ;
  signal N_28950_RETO_8 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_45\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_45\ : std_logic ;
  signal N_28951_RETO_0 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_46\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_46\ : std_logic ;
  signal N_28951_RETO_1 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_47\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_47\ : std_logic ;
  signal N_28951_RETO_2 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_48\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_48\ : std_logic ;
  signal N_28951_RETO_3 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_49\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_49\ : std_logic ;
  signal N_28951_RETO_4 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_50\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_50\ : std_logic ;
  signal N_28951_RETO_5 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_51\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_51\ : std_logic ;
  signal N_28951_RETO_6 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_52\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_52\ : std_logic ;
  signal N_28951_RETO_7 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_53\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_53\ : std_logic ;
  signal N_28951_RETO_8 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_54\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_54\ : std_logic ;
  signal N_28952_RETO_0 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_55\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_55\ : std_logic ;
  signal N_28952_RETO_1 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_56\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_56\ : std_logic ;
  signal N_28952_RETO_2 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_57\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_57\ : std_logic ;
  signal N_28952_RETO_3 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_58\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_58\ : std_logic ;
  signal N_28952_RETO_4 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_59\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_59\ : std_logic ;
  signal N_28952_RETO_5 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_60\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_60\ : std_logic ;
  signal N_28952_RETO_6 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_61\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_61\ : std_logic ;
  signal N_28952_RETO_7 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_62\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_62\ : std_logic ;
  signal N_28952_RETO_8 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_0\ : std_logic ;
  signal N_81248_0 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_1\ : std_logic ;
  signal N_81248_1 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506_1\ : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_4\ : std_logic ;
  signal N_81563_0 : std_logic ;
  signal \GRLFPC2_0.R.MK.RST_0\ : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_5\ : std_logic ;
  signal N_81563_1 : std_logic ;
  signal \GRLFPC2_0.R.MK.RST_1\ : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_6\ : std_logic ;
  signal N_81563_2 : std_logic ;
  signal \GRLFPC2_0.R.MK.RST_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3729_I_0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3729_I_0_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_5\ : std_logic ;
  signal N_32141_1_0 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10927_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_27_S_0_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10918_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0_0\ : std_logic ;
  signal N_55054_RETO_0 : std_logic ;
  signal \GRLFPC2_0.COMB.V.STATE0\ : std_logic ;
  signal \GRLFPC2_0.V.FSR.CEXC_0_SQMUXA0\ : std_logic ;
  signal \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA0\ : std_logic ;
  signal \GRLFPC2_0.V.FSR.CEXC_3_SQMUXA0\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0_1\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0_2\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0_3\ : std_logic ;
  signal \GRLFPC2_0.V.FSR.FTT_1_IV_I_A30\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN1_V.STATE0\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV0\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV0_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV0_1\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV0_2\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV0_3\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV0_4\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV0_5\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV0_6\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV0_7\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0_4\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0_5\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0_6\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0_7\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M20\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M20_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M20_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M20_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M20_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M20_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M20_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M20_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M20_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M30\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M30_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M300\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M300_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M30_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M30_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M30_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M30_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M30_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M30_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M30_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M300_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M300_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M300_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M300_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M300_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M300_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M300_7\ : std_logic ;
  signal N_2 : std_logic ;
  signal N_3 : std_logic ;
  signal N_4 : std_logic ;
  signal N_5 : std_logic ;
  signal N_6 : std_logic ;
  signal N_7 : std_logic ;
  signal N_8 : std_logic ;
  signal N_9 : std_logic ;
  signal N_10 : std_logic ;
  signal N_11 : std_logic ;
  signal N_12 : std_logic ;
  signal N_13 : std_logic ;
  signal N_14 : std_logic ;
  signal N_16 : std_logic ;
  signal N_17 : std_logic ;
  signal N_18 : std_logic ;
  signal N_19 : std_logic ;
  signal N_20 : std_logic ;
  signal N_21 : std_logic ;
  signal N_22 : std_logic ;
  signal N_23 : std_logic ;
  signal N_24 : std_logic ;
  signal N_25 : std_logic ;
  signal N_26 : std_logic ;
  signal N_27 : std_logic ;
  signal N_28 : std_logic ;
  signal N_29 : std_logic ;
  signal N_30 : std_logic ;
  signal N_31 : std_logic ;
  signal N_32 : std_logic ;
  signal N_33 : std_logic ;
  signal N_34 : std_logic ;
  signal N_35 : std_logic ;
  signal N_36 : std_logic ;
  signal N_37 : std_logic ;
  signal N_38 : std_logic ;
  signal N_39 : std_logic ;
  signal N_40 : std_logic ;
  signal N_41 : std_logic ;
  signal N_42 : std_logic ;
  signal N_43 : std_logic ;
  signal N_44 : std_logic ;
  signal N_45 : std_logic ;
  signal N_46 : std_logic ;
  signal N_47 : std_logic ;
  signal N_48 : std_logic ;
  signal N_49 : std_logic ;
  signal N_50 : std_logic ;
  signal N_51 : std_logic ;
  signal N_52 : std_logic ;
  signal N_53 : std_logic ;
  signal N_54 : std_logic ;
  signal N_55 : std_logic ;
  signal N_56 : std_logic ;
  signal N_57 : std_logic ;
  signal N_58 : std_logic ;
  signal N_59 : std_logic ;
  signal N_60 : std_logic ;
  signal N_61 : std_logic ;
  signal N_62 : std_logic ;
  signal N_63 : std_logic ;
  signal N_64 : std_logic ;
  signal N_65 : std_logic ;
  signal N_66 : std_logic ;
  signal N_67 : std_logic ;
  signal N_68 : std_logic ;
  signal N_69 : std_logic ;
  signal N_70 : std_logic ;
  signal N_71 : std_logic ;
  signal N_72 : std_logic ;
  signal N_73 : std_logic ;
  signal N_74 : std_logic ;
  signal N_75 : std_logic ;
  signal N_76 : std_logic ;
  signal N_77 : std_logic ;
  signal N_78 : std_logic ;
  signal N_79 : std_logic ;
  signal N_80 : std_logic ;
  signal N_81 : std_logic ;
  signal N_82 : std_logic ;
  signal N_83 : std_logic ;
  signal N_84 : std_logic ;
  signal N_85 : std_logic ;
  signal N_86 : std_logic ;
  signal N_87 : std_logic ;
  signal N_88 : std_logic ;
  signal N_89 : std_logic ;
  signal N_90 : std_logic ;
  signal N_91 : std_logic ;
  signal N_92 : std_logic ;
  signal N_93 : std_logic ;
  signal N_94 : std_logic ;
  signal N_95 : std_logic ;
  signal N_96 : std_logic ;
  signal N_97 : std_logic ;
  signal N_98 : std_logic ;
  signal N_99 : std_logic ;
  signal N_100 : std_logic ;
  signal N_101 : std_logic ;
  signal N_102 : std_logic ;
  signal N_103 : std_logic ;
  signal N_104 : std_logic ;
  signal N_105 : std_logic ;
  signal N_106 : std_logic ;
  signal N_107 : std_logic ;
  signal N_108 : std_logic ;
  signal N_109 : std_logic ;
  signal N_110 : std_logic ;
  signal N_111 : std_logic ;
  signal N_112 : std_logic ;
  signal N_113 : std_logic ;
  signal N_114 : std_logic ;
  signal N_115 : std_logic ;
  signal N_116 : std_logic ;
  signal N_117 : std_logic ;
  signal N_118 : std_logic ;
  signal N_119 : std_logic ;
  signal N_120 : std_logic ;
  signal N_121 : std_logic ;
  signal N_122 : std_logic ;
  signal N_123 : std_logic ;
  signal N_124 : std_logic ;
  signal N_125 : std_logic ;
  signal N_126 : std_logic ;
  signal N_127 : std_logic ;
  signal N_128 : std_logic ;
  signal N_129 : std_logic ;
  signal N_130 : std_logic ;
  signal N_131 : std_logic ;
  signal N_132 : std_logic ;
  signal N_133 : std_logic ;
  signal N_134 : std_logic ;
  signal N_135 : std_logic ;
  signal N_136 : std_logic ;
  signal N_137 : std_logic ;
  signal N_138 : std_logic ;
  signal N_139 : std_logic ;
  signal N_140 : std_logic ;
  signal N_141 : std_logic ;
  signal N_142 : std_logic ;
  signal N_143 : std_logic ;
  signal N_144 : std_logic ;
  signal N_145 : std_logic ;
  signal N_146 : std_logic ;
  signal N_147 : std_logic ;
  signal N_148 : std_logic ;
  signal N_149 : std_logic ;
  signal N_150 : std_logic ;
  signal N_151 : std_logic ;
  signal N_152 : std_logic ;
  signal N_153 : std_logic ;
  signal N_154 : std_logic ;
  signal N_155 : std_logic ;
  signal N_156 : std_logic ;
  signal N_157 : std_logic ;
  signal N_158 : std_logic ;
  signal N_159 : std_logic ;
  signal N_160 : std_logic ;
  signal N_161 : std_logic ;
  signal N_162 : std_logic ;
  signal N_163 : std_logic ;
  signal N_164 : std_logic ;
  signal N_165 : std_logic ;
  signal N_166 : std_logic ;
  signal N_167 : std_logic ;
  signal N_168 : std_logic ;
  signal N_169 : std_logic ;
  signal N_170 : std_logic ;
  signal N_171 : std_logic ;
  signal N_172 : std_logic ;
  signal N_173 : std_logic ;
  signal N_174 : std_logic ;
  signal N_175 : std_logic ;
  signal N_176 : std_logic ;
  signal N_177 : std_logic ;
  signal N_178 : std_logic ;
  signal N_179 : std_logic ;
  signal N_180 : std_logic ;
  signal N_181 : std_logic ;
  signal N_182 : std_logic ;
  signal N_183 : std_logic ;
  signal N_184 : std_logic ;
  signal N_185 : std_logic ;
  signal N_186 : std_logic ;
  signal N_187 : std_logic ;
  signal N_188 : std_logic ;
  signal N_189 : std_logic ;
  signal N_190 : std_logic ;
  signal N_191 : std_logic ;
  signal N_192 : std_logic ;
  signal N_193 : std_logic ;
  signal N_194 : std_logic ;
  signal N_195 : std_logic ;
  signal N_196 : std_logic ;
  signal N_197 : std_logic ;
  signal N_198 : std_logic ;
  signal N_199 : std_logic ;
  signal N_200 : std_logic ;
  signal N_201 : std_logic ;
  signal N_202 : std_logic ;
  signal N_203 : std_logic ;
  signal N_204 : std_logic ;
  signal N_205 : std_logic ;
  signal N_206 : std_logic ;
  signal N_207 : std_logic ;
  signal N_208 : std_logic ;
  signal N_209 : std_logic ;
  signal N_210 : std_logic ;
  signal N_211 : std_logic ;
  signal N_212 : std_logic ;
  signal N_213 : std_logic ;
  signal N_214 : std_logic ;
  signal N_215 : std_logic ;
  signal N_216 : std_logic ;
  signal N_217 : std_logic ;
  signal N_218 : std_logic ;
  signal N_219 : std_logic ;
  signal N_220 : std_logic ;
  signal N_221 : std_logic ;
  signal N_222 : std_logic ;
  signal N_223 : std_logic ;
  signal N_224 : std_logic ;
  signal N_225 : std_logic ;
  signal N_226 : std_logic ;
  signal N_227 : std_logic ;
  signal N_228 : std_logic ;
  signal N_229 : std_logic ;
  signal N_230 : std_logic ;
  signal N_231 : std_logic ;
  signal N_232 : std_logic ;
  signal N_233 : std_logic ;
  signal N_234 : std_logic ;
  signal N_235 : std_logic ;
  signal N_236 : std_logic ;
  signal N_237 : std_logic ;
  signal N_238 : std_logic ;
  signal N_239 : std_logic ;
  signal N_240 : std_logic ;
  signal N_241 : std_logic ;
  signal N_242 : std_logic ;
  signal N_243 : std_logic ;
  signal N_244 : std_logic ;
  signal N_245 : std_logic ;
  signal N_246 : std_logic ;
  signal N_247 : std_logic ;
  signal N_248 : std_logic ;
  signal N_249 : std_logic ;
  signal N_250 : std_logic ;
  signal N_251 : std_logic ;
  signal N_252 : std_logic ;
  signal N_253 : std_logic ;
  signal N_254 : std_logic ;
  signal N_255 : std_logic ;
  signal N_256 : std_logic ;
  signal N_257 : std_logic ;
  signal N_258 : std_logic ;
  signal N_259 : std_logic ;
  signal N_260 : std_logic ;
  signal N_261 : std_logic ;
  signal N_262 : std_logic ;
  signal N_263 : std_logic ;
  signal N_264 : std_logic ;
  signal N_265 : std_logic ;
  signal N_266 : std_logic ;
  signal N_267 : std_logic ;
  signal N_268 : std_logic ;
  signal N_269 : std_logic ;
  signal N_270 : std_logic ;
  signal N_271 : std_logic ;
  signal N_272 : std_logic ;
  signal N_273 : std_logic ;
  signal N_274 : std_logic ;
  signal N_275 : std_logic ;
  signal N_276 : std_logic ;
  signal N_277 : std_logic ;
  signal N_278 : std_logic ;
  signal N_279 : std_logic ;
  signal N_280 : std_logic ;
  signal N_281 : std_logic ;
  signal N_282 : std_logic ;
  signal N_283 : std_logic ;
  signal N_284 : std_logic ;
  signal N_285 : std_logic ;
  signal N_286 : std_logic ;
  signal N_287 : std_logic ;
  signal N_288 : std_logic ;
  signal N_289 : std_logic ;
  signal N_290 : std_logic ;
  signal N_291 : std_logic ;
  signal N_292 : std_logic ;
  signal N_293 : std_logic ;
  signal N_294 : std_logic ;
  signal N_295 : std_logic ;
  signal N_296 : std_logic ;
  signal N_297 : std_logic ;
  signal N_298 : std_logic ;
  signal N_299 : std_logic ;
  signal N_300 : std_logic ;
  signal N_301 : std_logic ;
  signal N_302 : std_logic ;
  signal N_303 : std_logic ;
  signal N_304 : std_logic ;
  signal N_305 : std_logic ;
  signal N_306 : std_logic ;
  signal N_307 : std_logic ;
  signal N_308 : std_logic ;
  signal N_309 : std_logic ;
  signal N_310 : std_logic ;
  signal N_311 : std_logic ;
  signal N_312 : std_logic ;
  signal N_313 : std_logic ;
  signal N_314 : std_logic ;
  signal N_315 : std_logic ;
  signal N_316 : std_logic ;
  signal N_317 : std_logic ;
  signal N_318 : std_logic ;
  signal N_319 : std_logic ;
  signal N_320 : std_logic ;
  signal N_321 : std_logic ;
  signal N_322 : std_logic ;
  signal N_323 : std_logic ;
  signal N_324 : std_logic ;
  signal N_325 : std_logic ;
  signal N_326 : std_logic ;
  signal N_327 : std_logic ;
  signal N_328 : std_logic ;
  signal N_329 : std_logic ;
  signal N_330 : std_logic ;
  signal N_331 : std_logic ;
  signal N_332 : std_logic ;
  signal N_333 : std_logic ;
  signal N_334 : std_logic ;
  signal N_335 : std_logic ;
  signal N_336 : std_logic ;
  signal N_337 : std_logic ;
  signal N_338 : std_logic ;
  signal N_339 : std_logic ;
  signal N_340 : std_logic ;
  signal N_341 : std_logic ;
  signal N_342 : std_logic ;
  signal N_343 : std_logic ;
  signal N_344 : std_logic ;
  signal N_345 : std_logic ;
  signal N_346 : std_logic ;
  signal N_347 : std_logic ;
  signal N_348 : std_logic ;
  signal N_349 : std_logic ;
  signal N_350 : std_logic ;
  signal N_351 : std_logic ;
  signal N_352 : std_logic ;
  signal N_353 : std_logic ;
  signal N_354 : std_logic ;
  signal N_355 : std_logic ;
  signal N_356 : std_logic ;
  signal N_357 : std_logic ;
  signal N_358 : std_logic ;
  signal N_359 : std_logic ;
  signal N_360 : std_logic ;
  signal N_361 : std_logic ;
  signal N_362 : std_logic ;
  signal N_363 : std_logic ;
  signal N_364 : std_logic ;
  signal N_365 : std_logic ;
  signal N_366 : std_logic ;
  signal N_367 : std_logic ;
  signal N_368 : std_logic ;
  signal N_369 : std_logic ;
  signal N_370 : std_logic ;
  signal N_371 : std_logic ;
  signal N_372 : std_logic ;
  signal N_373 : std_logic ;
  signal N_374 : std_logic ;
  signal N_375 : std_logic ;
  signal N_376 : std_logic ;
  signal N_377 : std_logic ;
  signal N_378 : std_logic ;
  signal N_379 : std_logic ;
  signal N_380 : std_logic ;
  signal N_381 : std_logic ;
  signal N_382 : std_logic ;
  signal N_383 : std_logic ;
  signal N_384 : std_logic ;
  signal N_385 : std_logic ;
  signal N_386 : std_logic ;
  signal N_387 : std_logic ;
  signal N_388 : std_logic ;
  signal N_389 : std_logic ;
  signal N_390 : std_logic ;
  signal N_391 : std_logic ;
  signal N_392 : std_logic ;
  signal N_393 : std_logic ;
  signal N_394 : std_logic ;
  signal N_395 : std_logic ;
  signal N_396 : std_logic ;
  signal N_397 : std_logic ;
  signal N_398 : std_logic ;
  signal N_399 : std_logic ;
  signal N_400 : std_logic ;
  signal N_401 : std_logic ;
  signal N_402 : std_logic ;
  signal N_403 : std_logic ;
  signal N_404 : std_logic ;
  signal N_405 : std_logic ;
  signal N_406 : std_logic ;
  signal N_407 : std_logic ;
  signal N_408 : std_logic ;
  signal N_409 : std_logic ;
  signal N_410 : std_logic ;
  signal N_411 : std_logic ;
  signal N_412 : std_logic ;
  signal N_413 : std_logic ;
  signal N_414 : std_logic ;
  signal N_415 : std_logic ;
  signal N_416 : std_logic ;
  signal N_417 : std_logic ;
  signal N_418 : std_logic ;
  signal N_419 : std_logic ;
  signal N_420 : std_logic ;
  signal N_421 : std_logic ;
  signal N_422 : std_logic ;
  signal N_423 : std_logic ;
  signal N_424 : std_logic ;
  signal N_425 : std_logic ;
  signal N_426 : std_logic ;
  signal N_427 : std_logic ;
  signal N_428 : std_logic ;
  signal N_429 : std_logic ;
  signal N_430 : std_logic ;
  signal N_431 : std_logic ;
  signal N_432 : std_logic ;
  signal N_433 : std_logic ;
  signal N_434 : std_logic ;
  signal N_0 : std_logic ;
  signal N_1_115 : std_logic ;
  signal N_2_116 : std_logic ;
  signal N_3_117 : std_logic ;
  signal N_4_118 : std_logic ;
  signal N_5_119 : std_logic ;
  signal N_6_120 : std_logic ;
  signal N_7_121 : std_logic ;
  signal N_8_122 : std_logic ;
  signal N_9_123 : std_logic ;
  signal N_10_124 : std_logic ;
  signal N_11_125 : std_logic ;
  signal N_12_126 : std_logic ;
  signal N_13_127 : std_logic ;
  signal N_14_128 : std_logic ;
  signal N_15_129 : std_logic ;
  signal N_16_130 : std_logic ;
  signal N_17_131 : std_logic ;
  signal N_18_132 : std_logic ;
  signal N_19_133 : std_logic ;
  signal N_20_134 : std_logic ;
  signal N_21_135 : std_logic ;
  signal N_22_136 : std_logic ;
  signal N_23_137 : std_logic ;
  signal N_24_138 : std_logic ;
  signal N_25_139 : std_logic ;
  signal N_26_140 : std_logic ;
  signal N_27_141 : std_logic ;
  signal N_28_142 : std_logic ;
  signal N_29_143 : std_logic ;
  signal N_30_144 : std_logic ;
  signal N_31_145 : std_logic ;
  signal N_32_146 : std_logic ;
  signal N_33_147 : std_logic ;
  signal N_34_148 : std_logic ;
  signal N_35_149 : std_logic ;
  signal N_36_150 : std_logic ;
  signal N_37_151 : std_logic ;
  signal N_38_152 : std_logic ;
  signal N_39_153 : std_logic ;
  signal N_40_154 : std_logic ;
  signal N_41_155 : std_logic ;
  signal N_42_156 : std_logic ;
  signal N_43_157 : std_logic ;
  signal N_44_158 : std_logic ;
  signal N_45_159 : std_logic ;
  signal N_46_160 : std_logic ;
  signal N_47_161 : std_logic ;
  signal N_48_162 : std_logic ;
  signal N_49_163 : std_logic ;
  signal N_50_164 : std_logic ;
  signal N_51_165 : std_logic ;
  signal N_52_166 : std_logic ;
  signal N_53_167 : std_logic ;
  signal N_54_168 : std_logic ;
  signal N_55_169 : std_logic ;
  signal N_56_170 : std_logic ;
  signal N_57_171 : std_logic ;
  signal N_58_172 : std_logic ;
  signal N_59_173 : std_logic ;
  signal N_60_174 : std_logic ;
  signal N_61_175 : std_logic ;
  signal N_62_176 : std_logic ;
  signal N_63_177 : std_logic ;
  signal N_64_178 : std_logic ;
  signal N_65_179 : std_logic ;
  signal N_66_180 : std_logic ;
  signal N_67_181 : std_logic ;
  signal N_68_182 : std_logic ;
  signal N_69_183 : std_logic ;
  signal N_70_184 : std_logic ;
  signal N_71_185 : std_logic ;
  signal N_72_186 : std_logic ;
  signal N_73_187 : std_logic ;
  signal N_74_188 : std_logic ;
  signal N_75_189 : std_logic ;
  signal N_76_190 : std_logic ;
  signal N_77_191 : std_logic ;
  signal N_78_192 : std_logic ;
  signal N_79_193 : std_logic ;
  signal N_80_194 : std_logic ;
  signal N_81_195 : std_logic ;
  signal N_82_196 : std_logic ;
  signal N_83_197 : std_logic ;
  signal N_84_198 : std_logic ;
  signal N_85_199 : std_logic ;
  signal N_86_200 : std_logic ;
  signal N_87_201 : std_logic ;
  signal N_88_202 : std_logic ;
  signal N_89_203 : std_logic ;
  signal N_90_204 : std_logic ;
  signal N_91_205 : std_logic ;
  signal N_92_206 : std_logic ;
  signal N_93_207 : std_logic ;
  signal N_94_208 : std_logic ;
  signal N_95_209 : std_logic ;
  signal N_96_210 : std_logic ;
  signal N_97_211 : std_logic ;
  signal N_98_212 : std_logic ;
  signal N_99_213 : std_logic ;
  signal N_100_214 : std_logic ;
  signal N_101_215 : std_logic ;
  signal N_102_216 : std_logic ;
  signal N_103_217 : std_logic ;
  signal N_104_218 : std_logic ;
  signal N_105_219 : std_logic ;
  signal N_106_220 : std_logic ;
  signal N_107_221 : std_logic ;
  signal N_108_222 : std_logic ;
  signal N_109_223 : std_logic ;
  signal N_110_224 : std_logic ;
  signal N_111_225 : std_logic ;
  signal N_112_226 : std_logic ;
  signal N_113_227 : std_logic ;
  signal N_114_228 : std_logic ;
  signal N_115_229 : std_logic ;
  signal N_116_230 : std_logic ;
  signal N_117_231 : std_logic ;
  signal N_118_232 : std_logic ;
  signal N_119_233 : std_logic ;
  signal N_120_234 : std_logic ;
  signal N_121_235 : std_logic ;
  signal N_122_236 : std_logic ;
  signal N_123_237 : std_logic ;
  signal N_124_238 : std_logic ;
  signal N_125_239 : std_logic ;
  signal N_126_240 : std_logic ;
  signal N_127_241 : std_logic ;
  signal N_128_242 : std_logic ;
  signal N_129_243 : std_logic ;
  signal N_130_244 : std_logic ;
  signal N_131_245 : std_logic ;
  signal N_132_246 : std_logic ;
  signal N_133_247 : std_logic ;
  signal N_134_248 : std_logic ;
  signal N_135_249 : std_logic ;
  signal N_136_250 : std_logic ;
  signal N_137_251 : std_logic ;
  signal N_138_252 : std_logic ;
  signal N_139_253 : std_logic ;
  signal N_140_254 : std_logic ;
  signal N_141_255 : std_logic ;
  signal N_142_256 : std_logic ;
  signal N_143_257 : std_logic ;
  signal N_144_258 : std_logic ;
  signal N_145_259 : std_logic ;
  signal N_146_260 : std_logic ;
  signal N_147_261 : std_logic ;
  signal N_148_262 : std_logic ;
  signal N_149_263 : std_logic ;
  signal N_150_264 : std_logic ;
  signal N_151_265 : std_logic ;
  signal N_152_266 : std_logic ;
  signal N_153_267 : std_logic ;
  signal N_154_268 : std_logic ;
  signal N_155_269 : std_logic ;
  signal N_156_270 : std_logic ;
  signal N_157_271 : std_logic ;
  signal N_158_272 : std_logic ;
  signal N_159_273 : std_logic ;
  signal N_160_274 : std_logic ;
  signal N_161_275 : std_logic ;
  signal N_162_276 : std_logic ;
  signal N_163_277 : std_logic ;
  signal N_599 : std_logic ;
  signal N_600 : std_logic ;
  signal N_601 : std_logic ;
  signal N_602 : std_logic ;
  signal N_603 : std_logic ;
  signal N_604 : std_logic ;
  signal N_605 : std_logic ;
  signal N_606 : std_logic ;
  signal N_607 : std_logic ;
  signal N_608 : std_logic ;
  signal N_609 : std_logic ;
  signal N_610 : std_logic ;
  signal N_611 : std_logic ;
  signal N_612 : std_logic ;
  signal N_613 : std_logic ;
  signal N_614 : std_logic ;
  signal N_615 : std_logic ;
  signal N_616 : std_logic ;
  signal N_617 : std_logic ;
  signal N_618 : std_logic ;
  signal N_619 : std_logic ;
  signal N_620 : std_logic ;
  signal N_621 : std_logic ;
  signal N_622 : std_logic ;
  signal N_623 : std_logic ;
  signal N_624 : std_logic ;
  signal N_625 : std_logic ;
  signal N_626 : std_logic ;
  signal N_627 : std_logic ;
  signal N_628 : std_logic ;
  signal N_629 : std_logic ;
  signal N_630 : std_logic ;
  signal N_631 : std_logic ;
  signal N_632 : std_logic ;
  signal N_633 : std_logic ;
  signal N_634 : std_logic ;
  signal N_635 : std_logic ;
  signal N_636 : std_logic ;
  signal N_637 : std_logic ;
  signal N_638 : std_logic ;
  signal N_639 : std_logic ;
  signal N_640 : std_logic ;
  signal N_641 : std_logic ;
  signal N_642 : std_logic ;
  signal N_643 : std_logic ;
  signal N_644 : std_logic ;
  signal N_645 : std_logic ;
  signal N_646 : std_logic ;
  signal N_647 : std_logic ;
  signal N_648 : std_logic ;
  signal N_649 : std_logic ;
  signal N_650 : std_logic ;
  signal N_651 : std_logic ;
  signal N_652 : std_logic ;
  signal N_653 : std_logic ;
  signal N_654 : std_logic ;
  signal N_655 : std_logic ;
  signal N_656 : std_logic ;
  signal N_657 : std_logic ;
  signal N_658 : std_logic ;
  signal N_659 : std_logic ;
  signal N_660 : std_logic ;
  signal N_661 : std_logic ;
  signal N_662 : std_logic ;
  signal N_663 : std_logic ;
  signal N_664 : std_logic ;
  signal N_665 : std_logic ;
  signal N_666 : std_logic ;
  signal N_667 : std_logic ;
  signal N_668 : std_logic ;
  signal N_669 : std_logic ;
  signal N_670 : std_logic ;
  signal N_671 : std_logic ;
  signal N_672 : std_logic ;
  signal N_673 : std_logic ;
  signal N_674 : std_logic ;
  signal N_675 : std_logic ;
  signal N_676 : std_logic ;
  signal N_677 : std_logic ;
  signal N_678 : std_logic ;
  signal N_679 : std_logic ;
  signal N_680 : std_logic ;
  signal N_681 : std_logic ;
  signal N_682 : std_logic ;
  signal N_683 : std_logic ;
  signal N_684 : std_logic ;
  signal N_685 : std_logic ;
  signal N_686 : std_logic ;
  signal N_687 : std_logic ;
  signal N_688 : std_logic ;
  signal N_689 : std_logic ;
  signal N_690 : std_logic ;
  signal N_691 : std_logic ;
  signal N_692 : std_logic ;
  signal N_693 : std_logic ;
  signal N_694 : std_logic ;
  signal N_695 : std_logic ;
  signal N_696 : std_logic ;
  signal N_697 : std_logic ;
  signal N_698 : std_logic ;
  signal N_699 : std_logic ;
  signal N_700 : std_logic ;
  signal N_701 : std_logic ;
  signal N_702 : std_logic ;
  signal N_703 : std_logic ;
  signal N_704 : std_logic ;
  signal N_705 : std_logic ;
  signal N_706 : std_logic ;
  signal N_707 : std_logic ;
  signal N_708 : std_logic ;
  signal N_709 : std_logic ;
  signal N_710 : std_logic ;
  signal N_711 : std_logic ;
  signal N_712 : std_logic ;
  signal N_713 : std_logic ;
  signal N_714 : std_logic ;
  signal N_715 : std_logic ;
  signal N_716 : std_logic ;
  signal N_717 : std_logic ;
  signal N_718 : std_logic ;
  signal N_719 : std_logic ;
  signal N_720 : std_logic ;
  signal N_721 : std_logic ;
  signal N_722 : std_logic ;
  signal N_723 : std_logic ;
  signal N_724 : std_logic ;
  signal N_725 : std_logic ;
  signal N_726 : std_logic ;
  signal CPO_EXCZ : std_logic ;
  signal CPO_CCVZ : std_logic ;
  signal CPO_LDLOCKZ : std_logic ;
  signal CPO_HOLDNZ : std_logic ;
  signal RFI1_REN1Z : std_logic ;
  signal RFI1_REN2Z : std_logic ;
  signal RFI1_WRENZ : std_logic ;
  signal RFI2_REN1Z : std_logic ;
  signal RFI2_REN2Z : std_logic ;
  signal RFI2_WRENZ : std_logic ;
begin
VCC <= '1';
GND <= '0';
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIE4D8_29_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"000000aa0000aa55")
port map (
sumout => N_26536,
cout => N_28672,
shareout => N_28673,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(29),
cin => GND,
sharein => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIJSIV_30_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000fcc00000c33c")
port map (
sumout => N_26538,
cout => N_28675,
shareout => N_28676,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(30),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(30),
cin => N_28672,
sharein => N_28673);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_RNIHPRK4_31_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_26540,
cout => N_28678,
shareout => N_28679,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(31),
cin => N_28675,
sharein => N_28676);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI8V4I9_32_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_26542,
cout => N_28681,
shareout => N_28682,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(32),
cin => N_28678,
sharein => N_28679);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIOANCJ_33_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_26544,
cout => N_28684,
shareout => N_28685,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(33),
cin => N_28681,
sharein => N_28682);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIQ1S171_34_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_26546,
cout => N_28687,
shareout => N_28688,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(34),
cin => N_28684,
sharein => N_28685);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI0G5CE2_35_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_26548,
cout => N_28690,
shareout => N_28691,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(35),
cin => N_28687,
sharein => N_28688);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIECO0T4_36_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_26550,
cout => N_28693,
shareout => N_28694,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(36),
cin => N_28690,
sharein => N_28691);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIC5U9Q9_37_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_26552,
cout => N_28696,
shareout => N_28697,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(37),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(37),
cin => N_28693,
sharein => N_28694);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIAN9SKJ_38_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_26554,
cout => N_28699,
shareout => N_28700,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(38),
cin => N_28696,
sharein => N_28697);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI8R01A71_39_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_26556,
cout => N_28702,
shareout => N_28703,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(39),
cin => N_28699,
sharein => N_28700);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIOAFAKE2_40_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_26558,
cout => N_28705,
shareout => N_28706,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(40),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(40),
cin => N_28702,
sharein => N_28703);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIQ9CT8T_41_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_26560,
cout => N_28708,
shareout => N_28709,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(41),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(41),
cin => N_28705,
sharein => N_28706);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI0863IQ1_42_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_26562,
cout => N_28711,
shareout => N_28712,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(42),
cin => N_28708,
sharein => N_28709);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIE4QE4L3_43_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_26564,
cout => N_28714,
shareout => N_28715,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(43),
cin => N_28711,
sharein => N_28712);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNICT169A3_44_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_26566,
cout => N_28717,
shareout => N_28718,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(44),
cin => N_28714,
sharein => N_28715);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIAFHKIK2_45_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_26568,
cout => N_28720,
shareout => N_28721,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(45),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(45),
cin => N_28717,
sharein => N_28718);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI8JGH591_46_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_26570,
cout => N_28723,
shareout => N_28724,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(46),
cin => N_28720,
sharein => N_28721);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI6REBBI2_47_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_26572,
cout => N_28726,
shareout => N_28727,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(47),
cin => N_28723,
sharein => N_28724);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI4BBVM41_48_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_26574,
cout => N_28729,
shareout => N_28730,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(48),
cin => N_28726,
sharein => N_28727);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI2B47E92_49_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_26576,
cout => N_28732,
shareout => N_28733,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(49),
cin => N_28729,
sharein => N_28730);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIIIMMSI_50_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_26578,
cout => N_28735,
shareout => N_28736,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(50),
cin => N_28732,
sharein => N_28733);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIK1RLP51_51_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_26580,
cout => N_28738,
shareout => N_28739,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(51),
cin => N_28735,
sharein => N_28736);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIQV3KJB2_52_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_26582,
cout => N_28741,
shareout => N_28742,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(52),
cin => N_28738,
sharein => N_28739);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI8SLG7N_53_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_26584,
cout => N_28744,
shareout => N_28745,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(53),
cin => N_28741,
sharein => N_28742);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI6LP9FE1_54_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_26586,
cout => N_28747,
shareout => N_28748,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(54),
cin => N_28744,
sharein => N_28745);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI471SUS2_55_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_26588,
cout => N_28750,
shareout => N_28751,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(55),
cin => N_28747,
sharein => N_28748);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI2BG0UP1_56_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_26590,
cout => N_28753,
shareout => N_28754,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(56),
cin => N_28750,
sharein => N_28751);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI0JE9SJ3_57_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_26592,
cout => N_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(57),
cin => N_28753,
sharein => N_28754);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIE4D8_0_29_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_26535,
cout => N_28759,
shareout => N_28760,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(29),
cin => GND,
sharein => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIUK7P_30_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_26537,
cout => N_28762,
shareout => N_28763,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(30),
cin => N_28759,
sharein => N_28760);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_RNI7A584_31_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_26539,
cout => N_28765,
shareout => N_28766,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(31),
cin => N_28762,
sharein => N_28763);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIK0OO8_32_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_26541,
cout => N_28768,
shareout => N_28769,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(32),
cin => N_28765,
sharein => N_28766);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIGDTPH_33_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_26543,
cout => N_28771,
shareout => N_28772,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(33),
cin => N_28768,
sharein => N_28769);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIA78S31_34_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_26545,
cout => N_28774,
shareout => N_28775,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(34),
cin => N_28771,
sharein => N_28772);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI0RT082_35_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_26547,
cout => N_28777,
shareout => N_28778,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(35),
cin => N_28774,
sharein => N_28775);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIE29AG4_36_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_26549,
cout => N_28780,
shareout => N_28781,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(36),
cin => N_28777,
sharein => N_28778);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNICHVS09_37_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_26551,
cout => N_28783,
shareout => N_28784,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(37),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(37),
cin => N_28780,
sharein => N_28781);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIAFC22I_38_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_26553,
cout => N_28786,
shareout => N_28787,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(38),
cin => N_28783,
sharein => N_28784);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI8B6D441_39_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_26555,
cout => N_28789,
shareout => N_28790,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(39),
cin => N_28786,
sharein => N_28787);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIOAQ2982_40_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_26557,
cout => N_28792,
shareout => N_28793,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(40),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(40),
cin => N_28789,
sharein => N_28790);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIQ92EIG_41_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_26559,
cout => N_28795,
shareout => N_28796,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(41),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(41),
cin => N_28792,
sharein => N_28793);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI08I4511_42_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_26561,
cout => N_28798,
shareout => N_28799,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(42),
cin => N_28795,
sharein => N_28796);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIE4IHA22_43_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_26563,
cout => N_28801,
shareout => N_28802,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(43),
cin => N_28798,
sharein => N_28799);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNICTHBL4_44_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_26565,
cout => N_28804,
shareout => N_28805,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(44),
cin => N_28801,
sharein => N_28802);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIAFHVA9_45_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_26567,
cout => N_28807,
shareout => N_28808,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(45),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(45),
cin => N_28804,
sharein => N_28805);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI8JG7MI_46_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_26569,
cout => N_28810,
shareout => N_28811,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(46),
cin => N_28807,
sharein => N_28808);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI6RENC51_47_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_26571,
cout => N_28813,
shareout => N_28814,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(47),
cin => N_28810,
sharein => N_28811);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI4BBNPA2_48_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_26573,
cout => N_28816,
shareout => N_28817,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(48),
cin => N_28813,
sharein => N_28814);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI2B4NJL_49_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_26575,
cout => N_28819,
shareout => N_28820,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(49),
cin => N_28816,
sharein => N_28817);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIIIMM7B1_50_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_26577,
cout => N_28822,
shareout => N_28823,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(50),
cin => N_28819,
sharein => N_28820);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIK1RLFM2_51_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_26579,
cout => N_28825,
shareout => N_28826,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(51),
cin => N_28822,
sharein => N_28823);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIQV3KVC1_52_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_26581,
cout => N_28828,
shareout => N_28829,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(52),
cin => N_28825,
sharein => N_28826);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI8SLGVP2_53_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_26583,
cout => N_28831,
shareout => N_28832,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(53),
cin => N_28828,
sharein => N_28829);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI6LP9VJ1_54_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_26585,
cout => N_28834,
shareout => N_28835,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(54),
cin => N_28831,
sharein => N_28832);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI471SU73_55_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_26587,
cout => N_28837,
shareout => N_28838,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(55),
cin => N_28834,
sharein => N_28835);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI2BG0UF2_56_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_26589,
cout => N_28840,
shareout => N_28841,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(56),
cin => N_28837,
sharein => N_28838);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI0JE9SV_57_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_26591,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(57),
cin => N_28840,
sharein => N_28841);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN8_TEMP_U_RNIS4RU_0_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000ee8800009966")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(0),
cout => N_28846,
shareout => N_28847,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5410\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10560\,
cin => GND,
sharein => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI5JCG3_1_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(1),
cout => N_28849,
shareout => N_28850,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5391\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(1),
cin => N_28846,
sharein => N_28847);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIO5A67_2_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(2),
cout => N_28852,
shareout => N_28853,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(2),
cin => N_28849,
sharein => N_28850);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI0J5IE_3_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(3),
cout => N_28855,
shareout => N_28856,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(3),
cin => N_28852,
sharein => N_28853);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIILS9T_4_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(4),
cout => N_28858,
shareout => N_28859,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(4),
cin => N_28855,
sharein => N_28856);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIO2BPQ1_5_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(5),
cout => N_28861,
shareout => N_28862,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(5),
cin => N_28858,
sharein => N_28859);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI658OL3_6_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(6),
cout => N_28864,
shareout => N_28865,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(6),
cin => N_28861,
sharein => N_28862);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI4I2MB7_7_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(7),
cout => N_28867,
shareout => N_28868,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(7),
cin => N_28864,
sharein => N_28865);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI2KNHNE_8_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(8),
cout => N_28870,
shareout => N_28871,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(8),
cin => N_28867,
sharein => N_28868);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI0029FT_9_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(9),
cout => N_28873,
shareout => N_28874,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(9),
cin => N_28870,
sharein => N_28871);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIMRGQUQ1_10_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(10),
cout => N_28876,
shareout => N_28877,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(10),
cin => N_28873,
sharein => N_28874);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI4JETTL3_11_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(11),
cout => N_28879,
shareout => N_28880,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(11),
cin => N_28876,
sharein => N_28877);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI22A3SB3_12_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(12),
cout => N_28882,
shareout => N_28883,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(12),
cin => N_28879,
sharein => N_28880);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI001FON2_13_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(13),
cout => N_28885,
shareout => N_28886,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(13),
cin => N_28882,
sharein => N_28883);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIURE6HF1_14_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(14),
cout => N_28888,
shareout => N_28889,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(14),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(14),
cin => N_28885,
sharein => N_28886);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNISJAL2V2_15_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(15),
cout => N_28891,
shareout => N_28892,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(15),
cin => N_28888,
sharein => N_28889);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIQ32J5U1_16_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(16),
cout => N_28894,
shareout => N_28895,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(16),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(16),
cin => N_28891,
sharein => N_28892);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIO3HEBS3_17_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(17),
cout => N_28897,
shareout => N_28898,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(17),
cin => N_28894,
sharein => N_28895);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIM3F5NO3_18_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(18),
cout => N_28900,
shareout => N_28901,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(18),
cin => N_28897,
sharein => N_28898);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIK3BJEH3_19_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(19),
cout => N_28903,
shareout => N_28904,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(19),
cin => N_28900,
sharein => N_28901);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI4B3FT23_20_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(20),
cout => N_28906,
shareout => N_28907,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(20),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(20),
cin => N_28903,
sharein => N_28904);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI6QJ6R52_21_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(21),
cout => N_28909,
shareout => N_28910,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(21),
cin => N_28906,
sharein => N_28907);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNICOKLMB_22_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(22),
cout => N_28912,
shareout => N_28913,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(22),
cin => N_28909,
sharein => N_28910);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIQKMJDN_23_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(23),
cout => N_28915,
shareout => N_28916,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(23),
cin => N_28912,
sharein => N_28913);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIODQFRE1_24_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(24),
cout => N_28918,
shareout => N_28919,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(24),
cin => N_28915,
sharein => N_28916);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIMV18NT2_25_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(25),
cout => N_28921,
shareout => N_28922,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(25),
cin => N_28918,
sharein => N_28919);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIK3HOER1_26_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(26),
cout => N_28924,
shareout => N_28925,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(26),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(26),
cin => N_28921,
sharein => N_28922);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIIBFPTM3_27_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(27),
cout => N_28927,
shareout => N_28928,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(27),
cin => N_28924,
sharein => N_28925);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIGRBRRD3_28_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(28),
cout => N_28930,
shareout => N_28931,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(28),
cin => N_28927,
sharein => N_28928);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI0NNMNR2_28_\: stratixii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000000000000000")
port map (
sumout => N_26534,
cout => N_3,
cin => N_28930,
sharein => N_28931);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_21_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_22\(35),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21.Z_CARRY_0\,
dataf => N_57572,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(333),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57566);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_21_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_79\(34),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21.Z_CARRY_1\,
dataf => N_57578,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_21\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_21_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_136\(33),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21.Z_CARRY_2\,
dataf => N_57579,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_78\(35),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_21_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(21),
cout => N_57564,
dataf => N_57587,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_135\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_20_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_21\(36),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20.Z_CARRY_0\,
dataf => N_57595,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(332),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57562);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_20_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_78\(35),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20.Z_CARRY_1\,
dataf => N_57601,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_20\(37),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_20_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_135\(34),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20.Z_CARRY_2\,
dataf => N_57602,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_77\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_20_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(20),
cout => N_57560,
dataf => N_57610,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_134\(35),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_19_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_20\(37),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19.Z_CARRY_0\,
dataf => N_57618,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(331),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57558);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_19_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_77\(36),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19.Z_CARRY_1\,
dataf => N_57624,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_19\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_19_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_134\(35),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19.Z_CARRY_2\,
dataf => N_57625,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_76\(37),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_19_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(19),
cout => N_57556,
dataf => N_57633,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_133\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_18_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_19\(38),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18.Z_CARRY_0\,
dataf => N_57641,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(330),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57554);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_18_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_76\(37),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18.Z_CARRY_1\,
dataf => N_57647,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_18\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_18_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_133\(36),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18.Z_CARRY_2\,
dataf => N_57648,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_75\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_18_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(18),
cout => N_57552,
dataf => N_57656,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_132\(37),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_17_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_18\(39),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17.Z_CARRY_0\,
dataf => N_57664,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(329),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57550);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_17_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_75\(38),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17.Z_CARRY_1\,
dataf => N_57670,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_17\(40),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_17_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_132\(37),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17.Z_CARRY_2\,
dataf => N_57671,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_74\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_17_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(17),
cout => N_57548,
dataf => N_57679,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_131\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_16_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_17\(40),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16.Z_CARRY_0\,
dataf => N_57687,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(328),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57546);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_16_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_74\(39),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16.Z_CARRY_1\,
dataf => N_57693,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_16\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_16_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_131\(38),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16.Z_CARRY_2\,
dataf => N_57694,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_73\(40),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_16_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(16),
cout => N_57544,
dataf => N_57702,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_130\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_15_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_16\(41),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15.Z_CARRY_0\,
dataf => N_57710,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(327),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57542);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_15_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_73\(40),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15.Z_CARRY_1\,
dataf => N_57716,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_15\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_15_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_130\(39),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15.Z_CARRY_2\,
dataf => N_57717,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_72\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_15_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(15),
cout => N_57540,
dataf => N_57725,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_129\(40),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_14_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_15\(42),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14.Z_CARRY_0\,
dataf => N_57733,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(326),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57538);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_14_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_72\(41),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14.Z_CARRY_1\,
dataf => N_57739,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_14\(43),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_14_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_129\(40),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14.Z_CARRY_2\,
dataf => N_57740,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_71\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_14_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(14),
cout => N_57536,
dataf => N_57748,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_128\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_13_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_14\(43),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13.Z_CARRY_0\,
dataf => N_57756,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(325),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57534);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_13_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_71\(42),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13.Z_CARRY_1\,
dataf => N_57762,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_13\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_13_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_128\(41),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13.Z_CARRY_2\,
dataf => N_57763,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_70\(43),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_13_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(13),
cout => N_57532,
dataf => N_57771,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_127\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_12_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_13\(44),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12.Z_CARRY_0\,
dataf => N_57779,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(324),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57530);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_12_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_70\(43),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12.Z_CARRY_1\,
dataf => N_57785,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_12\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_12_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_127\(42),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12.Z_CARRY_2\,
dataf => N_57786,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_69\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_12_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(12),
cout => N_57528,
dataf => N_57794,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_126\(43),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_11_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_12\(45),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11.Z_CARRY_0\,
dataf => N_57802,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(323),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57526);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_11_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_69\(44),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11.Z_CARRY_1\,
dataf => N_57808,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_11\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_11_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_126\(43),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11.Z_CARRY_2\,
dataf => N_57809,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_68\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_11_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(11),
cout => N_57524,
dataf => N_57817,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_125\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_10_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_11\(46),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10.Z_CARRY_0\,
dataf => N_57825,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(322),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57522);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_10_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_68\(45),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10.Z_CARRY_1\,
dataf => N_57831,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_10\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_10_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_125\(44),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10.Z_CARRY_2\,
dataf => N_57832,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_67\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_10_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(10),
cout => N_57520,
dataf => N_57840,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_124\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_9_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_10\(47),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9.Z_CARRY_0\,
dataf => N_57848,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(321),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57518);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_9_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_67\(46),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9.Z_CARRY_1\,
dataf => N_57854,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_9\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_9_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_124\(45),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9.Z_CARRY_2\,
dataf => N_57855,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_66\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_9_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(9),
cout => N_57516,
dataf => N_57863,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_123\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_8_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_9\(48),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8.Z_CARRY_0\,
dataf => N_57871,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(320),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57514);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_8_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_66\(47),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8.Z_CARRY_1\,
dataf => N_57877,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_8\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_8_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_123\(46),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8.Z_CARRY_2\,
dataf => N_57878,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_65\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_8_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(8),
cout => N_57512,
dataf => N_57886,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_122\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_36_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_37\(20),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36.Z_CARRY_0\,
dataf => N_57894,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(348),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_57510);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_36_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_94\(19),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36.Z_CARRY_1\,
dataf => N_57900,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_36\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_36_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_151\(18),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36.Z_CARRY_2\,
dataf => N_57901,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_93\(20),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_36_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(36),
cout => N_57508,
dataf => N_57909,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_150\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_35_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_36\(21),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35.Z_CARRY_0\,
dataf => N_57917,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(347),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_57506);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_35_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_93\(20),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35.Z_CARRY_1\,
dataf => N_57923,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_35\(22),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_35_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_150\(19),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35.Z_CARRY_2\,
dataf => N_57924,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_92\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_35_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(35),
cout => N_57504,
dataf => N_57932,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_149\(20),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_34_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_35\(22),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34.Z_CARRY_0\,
dataf => N_57940,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(346),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_57502);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_34_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_92\(21),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34.Z_CARRY_1\,
dataf => N_57946,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_34\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_34_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_149\(20),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34.Z_CARRY_2\,
dataf => N_57947,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_91\(22),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_34_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(34),
cout => N_57500,
dataf => N_57955,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_148\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_33_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_34\(23),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33.Z_CARRY_0\,
dataf => N_57963,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(345),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57498);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_33_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_91\(22),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33.Z_CARRY_1\,
dataf => N_57969,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_33\(24),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_33_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_148\(21),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33.Z_CARRY_2\,
dataf => N_57970,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_90\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_33_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(33),
cout => N_57496,
dataf => N_57978,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_147\(22),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_32_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_33\(24),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32.Z_CARRY_0\,
dataf => N_57986,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(344),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57494);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_32_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_90\(23),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32.Z_CARRY_1\,
dataf => N_57992,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_32\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_32_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_147\(22),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32.Z_CARRY_2\,
dataf => N_57993,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_89\(24),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_32_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(32),
cout => N_57492,
dataf => N_58001,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_146\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_31_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_32\(25),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31.Z_CARRY_0\,
dataf => N_58009,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(343),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57490);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_31_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_89\(24),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31.Z_CARRY_1\,
dataf => N_58015,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_31\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_31_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_146\(23),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31.Z_CARRY_2\,
dataf => N_58016,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_88\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_31_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(31),
cout => N_57488,
dataf => N_58024,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_145\(24),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_30_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_31\(26),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30.Z_CARRY_0\,
dataf => N_58032,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(342),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57486);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_30_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_88\(25),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30.Z_CARRY_1\,
dataf => N_58038,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_30\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_30_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_145\(24),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30.Z_CARRY_2\,
dataf => N_58039,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_87\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_30_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(30),
cout => N_57484,
dataf => N_58047,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_144\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_29_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_30\(27),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29.Z_CARRY_0\,
dataf => N_58055,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(341),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57482);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_29_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_87\(26),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29.Z_CARRY_1\,
dataf => N_58061,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_29\(28),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_29_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_144\(25),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29.Z_CARRY_2\,
dataf => N_58062,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_86\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_29_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(29),
cout => N_57480,
dataf => N_58070,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_143\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_28_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_29\(28),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28.Z_CARRY_0\,
dataf => N_58078,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(340),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57478);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_28_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_86\(27),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28.Z_CARRY_1\,
dataf => N_58084,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_28\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_28_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_143\(26),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28.Z_CARRY_2\,
dataf => N_58085,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_85\(28),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_28_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(28),
cout => N_57476,
dataf => N_58093,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_142\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_27_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_28\(29),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27.Z_CARRY_0\,
dataf => N_58101,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(339),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57474);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_27_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_85\(28),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27.Z_CARRY_1\,
dataf => N_58107,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_27\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_27_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_142\(27),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27.Z_CARRY_2\,
dataf => N_58108,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_84\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_27_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(27),
cout => N_57472,
dataf => N_58116,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_141\(28),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_26_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_27\(30),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26.Z_CARRY_0\,
dataf => N_58124,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(338),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57470);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_26_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_84\(29),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26.Z_CARRY_1\,
dataf => N_58130,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_26\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_26_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_141\(28),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26.Z_CARRY_2\,
dataf => N_58131,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_83\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_26_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(26),
cout => N_57468,
dataf => N_58139,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_140\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_25_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_26\(31),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25.Z_CARRY_0\,
dataf => N_58147,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(337),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57466);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_25_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_83\(30),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25.Z_CARRY_1\,
dataf => N_58153,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_25\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_25_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_140\(29),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25.Z_CARRY_2\,
dataf => N_58154,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_82\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_25_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(25),
cout => N_57464,
dataf => N_58162,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_139\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_24_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_25\(32),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24.Z_CARRY_0\,
dataf => N_58170,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(336),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57462);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_24_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_82\(31),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24.Z_CARRY_1\,
dataf => N_58176,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_24\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_24_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_139\(30),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24.Z_CARRY_2\,
dataf => N_58177,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_81\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_24_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(24),
cout => N_57460,
dataf => N_58185,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_138\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_23_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_24\(33),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23.Z_CARRY_0\,
dataf => N_58193,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(335),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57458);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_23_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_81\(32),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23.Z_CARRY_1\,
dataf => N_58199,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_23\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_23_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_138\(31),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23.Z_CARRY_2\,
dataf => N_58200,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_80\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_23_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(23),
cout => N_57456,
dataf => N_58208,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_137\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_22_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_23\(34),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22.Z_CARRY_0\,
dataf => N_58216,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(334),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57454);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_22_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_80\(33),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22.Z_CARRY_1\,
dataf => N_58222,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_22\(35),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_22_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_137\(32),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22.Z_CARRY_2\,
dataf => N_58223,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_79\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_22_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(22),
cout => N_57452,
dataf => N_58231,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_136\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_51_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_52\(5),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51.Z_CARRY_0\,
dataf => N_58239,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(363),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_57450);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_51_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_109\(4),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51.Z_CARRY_1\,
dataf => N_58245,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_51\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_51_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_166\(3),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51.Z_CARRY_2\,
dataf => N_58246,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_108\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_51_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(51),
cout => N_57448,
dataf => N_58254,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_165\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_50_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_51\(6),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50.Z_CARRY_0\,
dataf => N_58262,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(362),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_57446);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_50_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_108\(5),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50.Z_CARRY_1\,
dataf => N_58268,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_50\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_50_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_165\(4),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50.Z_CARRY_2\,
dataf => N_58269,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_107\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_50_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(50),
cout => N_57444,
dataf => N_58277,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_164\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_49_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_50\(7),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49.Z_CARRY_0\,
dataf => N_58285,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(361),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_57442);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_49_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_107\(6),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49.Z_CARRY_1\,
dataf => N_58291,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_49\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_49_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_164\(5),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49.Z_CARRY_2\,
dataf => N_58292,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_106\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_49_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(49),
cout => N_57440,
dataf => N_58300,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_163\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_48_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_49\(8),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48.Z_CARRY_0\,
dataf => N_58308,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(360),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_57438);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_48_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_106\(7),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48.Z_CARRY_1\,
dataf => N_58314,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_48\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_48_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_163\(6),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48.Z_CARRY_2\,
dataf => N_58315,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_105\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_48_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(48),
cout => N_57436,
dataf => N_58323,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_162\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_47_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_48\(9),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47.Z_CARRY_0\,
dataf => N_58331,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(359),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_57434);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_47_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_105\(8),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47.Z_CARRY_1\,
dataf => N_58337,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_47\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_47_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_162\(7),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47.Z_CARRY_2\,
dataf => N_58338,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_104\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_47_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(47),
cout => N_57432,
dataf => N_58346,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_161\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_46_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_47\(10),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46.Z_CARRY_0\,
dataf => N_58354,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(358),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_57430);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_46_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_104\(9),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46.Z_CARRY_1\,
dataf => N_58360,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_46\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_46_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_161\(8),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46.Z_CARRY_2\,
dataf => N_58361,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_103\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_46_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(46),
cout => N_57428,
dataf => N_58369,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_160\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_45_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_46\(11),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45.Z_CARRY_0\,
dataf => N_58377,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(357),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_57426);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_45_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_103\(10),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45.Z_CARRY_1\,
dataf => N_58383,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_45\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_45_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_160\(9),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45.Z_CARRY_2\,
dataf => N_58384,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_102\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_45_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(45),
cout => N_57424,
dataf => N_58392,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_159\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_44_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_45\(12),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44.Z_CARRY_0\,
dataf => N_58400,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(356),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_57422);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_44_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_102\(11),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44.Z_CARRY_1\,
dataf => N_58406,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_44\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_44_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_159\(10),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44.Z_CARRY_2\,
dataf => N_58407,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_101\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_44_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(44),
cout => N_57420,
dataf => N_58415,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_158\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_43_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_44\(13),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43.Z_CARRY_0\,
dataf => N_58423,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(355),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_57418);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_43_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_101\(12),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43.Z_CARRY_1\,
dataf => N_58429,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_43\(14),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_43_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_158\(11),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43.Z_CARRY_2\,
dataf => N_58430,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_100\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_43_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(43),
cout => N_57416,
dataf => N_58438,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_157\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_42_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_43\(14),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42.Z_CARRY_0\,
dataf => N_58446,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(354),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_57414);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_42_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_100\(13),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42.Z_CARRY_1\,
dataf => N_58452,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_42\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_42_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_157\(12),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42.Z_CARRY_2\,
dataf => N_58453,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_99\(14),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_42_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(42),
cout => N_57412,
dataf => N_58461,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_156\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_41_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_42\(15),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41.Z_CARRY_0\,
dataf => N_58469,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(353),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_57410);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_41_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_99\(14),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41.Z_CARRY_1\,
dataf => N_58475,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_41\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_41_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_156\(13),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41.Z_CARRY_2\,
dataf => N_58476,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_98\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_41_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(41),
cout => N_57408,
dataf => N_58484,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_155\(14),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_40_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_41\(16),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40.Z_CARRY_0\,
dataf => N_58492,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(352),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_57406);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_40_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_98\(15),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40.Z_CARRY_1\,
dataf => N_58498,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_40\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_40_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_155\(14),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40.Z_CARRY_2\,
dataf => N_58499,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_97\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_40_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(40),
cout => N_57404,
dataf => N_58507,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_154\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_39_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_40\(17),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39.Z_CARRY_0\,
dataf => N_58515,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(351),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_57402);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_39_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_97\(16),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39.Z_CARRY_1\,
dataf => N_58521,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_39\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_39_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_154\(15),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39.Z_CARRY_2\,
dataf => N_58522,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_96\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_39_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(39),
cout => N_57400,
dataf => N_58530,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_153\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_38_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_39\(18),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38.Z_CARRY_0\,
dataf => N_58538,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(350),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_57398);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_38_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_96\(17),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38.Z_CARRY_1\,
dataf => N_58544,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_38\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_38_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_153\(16),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38.Z_CARRY_2\,
dataf => N_58545,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_95\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_38_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(38),
cout => N_57396,
dataf => N_58553,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_152\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_37_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_38\(19),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37.Z_CARRY_0\,
dataf => N_58561,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(349),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_57394);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_37_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_95\(18),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37.Z_CARRY_1\,
dataf => N_58567,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_37\(20),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_37_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_152\(17),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37.Z_CARRY_2\,
dataf => N_58568,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_94\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_37_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(37),
cout => N_57392,
dataf => N_58576,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_151\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff000000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(0),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(257),
cin => N_81973);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff000000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(1),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(243),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(256),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff000000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(2),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(255),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff000000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(3),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(241),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(254),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CARRY_4: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff000000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(4),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(240),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(253),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CARRY_5: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff000000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(5),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(239),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(252),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_4\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CARRY_6: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff000000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(6),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(238),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(251),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_5\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CARRY_7: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff000000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(7),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(237),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(250),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_6\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CARRY_8: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff000000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(8),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(249),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_7\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CARRY_9: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff000000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(9),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_9\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(248),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_8\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CARRY_10: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff000000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(10),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_10\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(247),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_9\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CARRY_11: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff000000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(11),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_11\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_10\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CARRY_12: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff000000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(12),
cout => N_4,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(232),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(245),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_11\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_7_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_8\(49),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7.Z_CARRY_0\,
dataf => N_58586,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(319),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57388);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_7_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_65\(48),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7.Z_CARRY_1\,
dataf => N_58592,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_7\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_7_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_122\(47),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7.Z_CARRY_2\,
dataf => N_58593,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_64\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_7_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(7),
cout => N_57386,
dataf => N_58601,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_121\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_6_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_7\(50),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6.Z_CARRY_0\,
dataf => N_58609,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(318),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57384);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_6_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_64\(49),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6.Z_CARRY_1\,
dataf => N_58615,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_6\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_6_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_121\(48),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6.Z_CARRY_2\,
dataf => N_58616,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_63\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_6_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(6),
cout => N_57382,
dataf => N_58624,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_120\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_5_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_6\(51),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5.Z_CARRY_0\,
dataf => N_58632,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(317),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57380);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_5_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_63\(50),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5.Z_CARRY_1\,
dataf => N_58638,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_5\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_5_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_120\(49),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5.Z_CARRY_2\,
dataf => N_58639,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_62\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_5_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(5),
cout => N_57378,
dataf => N_58647,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_119\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_4_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_5\(52),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4.Z_CARRY_0\,
dataf => N_58657,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(316),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_57376);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_4_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000ff0")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_62\(51),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4.Z_CARRY_1\,
dataf => N_58667,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_12239\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5771\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_4_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000ff0")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_119\(50),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4.Z_CARRY_2\,
dataf => N_58668,
datad => N_34177,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6583\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_4_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000ff0")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(4),
cout => N_57374,
dataf => N_58672,
datad => N_58671,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_60.Z_1_CO0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6961\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_55_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_56\(1),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55.Z_CARRY_0\,
dataf => N_58677,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(367),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_57372);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_55_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_113\(0),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55.Z_CARRY_1\,
dataf => N_58683,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_55\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_55_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SCLSBS_1\(1),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55.Z_CARRY_2\,
dataf => N_58684,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_112\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_55_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000c00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(55),
cout => N_57370,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI\(0),
datad => N_58692,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_54_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_55\(2),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54.Z_CARRY_0\,
dataf => N_58700,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(366),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_57368);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_54_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_112\(1),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54.Z_CARRY_1\,
dataf => N_58706,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_54\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_54_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI\(0),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54.Z_CARRY_2\,
dataf => N_58707,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_111\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_54_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(54),
cout => N_57366,
dataf => N_58715,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_168\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_53_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_54\(3),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53.Z_CARRY_0\,
dataf => N_58723,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(365),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_57364);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_53_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_111\(2),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53.Z_CARRY_1\,
dataf => N_58729,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_53\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_53_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_168\(1),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53.Z_CARRY_2\,
dataf => N_58730,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_110\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_53_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(53),
cout => N_57362,
dataf => N_58738,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_167\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_52_Z_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_53\(4),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52.Z_CARRY_0\,
dataf => N_58746,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(364),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_57360);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_52_Z_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_110\(3),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52.Z_CARRY_1\,
dataf => N_58752,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_52\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_52_Z_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_167\(2),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52.Z_CARRY_2\,
dataf => N_58753,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_109\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_52_Z_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(52),
cout => N_57358,
dataf => N_58761,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_166\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff0000f0cc")
port map (
sumout => \GRLFPC2_0.FPO.EXP\(0),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10878\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10865\,
cin => N_57356);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff0000f3c0")
port map (
sumout => \GRLFPC2_0.FPO.EXP\(1),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10866\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10879\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff0000f3c0")
port map (
sumout => \GRLFPC2_0.FPO.EXP\(2),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10867\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10880\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff0000f3c0")
port map (
sumout => \GRLFPC2_0.FPO.EXP\(3),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10868\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10881\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_4: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff0000f3c0")
port map (
sumout => \GRLFPC2_0.FPO.EXP\(4),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10869\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10882\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_5: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff0000fc30")
port map (
sumout => \GRLFPC2_0.FPO.EXP\(5),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10883\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10870\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_4\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_6: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff0000fc30")
port map (
sumout => \GRLFPC2_0.FPO.EXP\(6),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10884\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10870\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_5\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_7: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff0000fc30")
port map (
sumout => \GRLFPC2_0.FPO.EXP\(7),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10885\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10872\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_6\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_8: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff0000fc30")
port map (
sumout => \GRLFPC2_0.FPO.EXP\(8),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10886\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10872\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_7\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_9: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff0000f3c0")
port map (
sumout => \GRLFPC2_0.FPO.EXP\(9),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_9\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10872\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10887\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_8\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_10: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cc330000f000")
port map (
sumout => \GRLFPC2_0.FPO.EXP\(10),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_10\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5301\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10888\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_9\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_11: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cc330000f000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\(11),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_11\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5343\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10889\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_10\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_12: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cc330000f000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\(12),
cout => N_5,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5339\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10890\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_11\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_3_0_RNIQC7P: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ccff0000f000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_57\(0),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(368),
datad => N_58821,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
cin => N_57354);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_0_RNI5BMN1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00003000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SBLSBS_1\(1),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_56\(1),
datad => N_58827,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_1_0_RNI8AOM3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SCLSBS_2\(0),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_2\,
dataf => N_58828,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_113\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_1_0_RNI8AOM3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_954\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_3\,
dataf => VCC,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_1_0_RNIOCGF7: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN25_NOTPROP\,
cout => N_57352,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SCLSBS_1\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_1_0_RNIOCGF7_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_4\,
cout => N_6,
cin => N_57352);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_RNITKAC_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57354,
datad => N_58820,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000f0cc")
port map (
cout => N_57356,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(35),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_52_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(109),
cin => N_57358);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_52_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57360,
datad => N_58745,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_53_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(110),
cin => N_57362);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_53_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57364,
datad => N_58722,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_54_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(111),
cin => N_57366);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_54_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57368,
datad => N_58699,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_55_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(112),
cin => N_57370);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_55_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57372,
datad => N_58676,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_4_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(61),
cin => N_57374);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_4_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57376,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10634\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_5_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(62),
cin => N_57378);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_5_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57380,
datad => N_58631,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_6_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(63),
cin => N_57382);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_6_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57384,
datad => N_58608,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_7_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(64),
cin => N_57386);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_7_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57388,
datad => N_58585,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_37_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(94),
cin => N_57392);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_37_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57394,
datad => N_58560,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_38_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(95),
cin => N_57396);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_38_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57398,
datad => N_58537,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_39_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(96),
cin => N_57400);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_39_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57402,
datad => N_58514,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_40_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(97),
cin => N_57404);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_40_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57406,
datad => N_58491,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_41_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(98),
cin => N_57408);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_41_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57410,
datad => N_58468,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_42_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(99),
cin => N_57412);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_42_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57414,
datad => N_58445,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_43_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(100),
cin => N_57416);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_43_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57418,
datad => N_58422,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_44_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(101),
cin => N_57420);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_44_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57422,
datad => N_58399,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_45_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(102),
cin => N_57424);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_45_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57426,
datad => N_58376,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_46_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(103),
cin => N_57428);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_46_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57430,
datad => N_58353,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_47_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(104),
cin => N_57432);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_47_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57434,
datad => N_58330,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_48_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(105),
cin => N_57436);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_48_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57438,
datad => N_58307,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_49_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(106),
cin => N_57440);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_49_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57442,
datad => N_58284,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_50_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(107),
cin => N_57444);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_50_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57446,
datad => N_58261,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_51_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(108),
cin => N_57448);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_51_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57450,
datad => N_58238,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_22_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(79),
cin => N_57452);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_22_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57454,
datad => N_58215,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_23_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(80),
cin => N_57456);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_23_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57458,
datad => N_58192,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_24_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(81),
cin => N_57460);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_24_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57462,
datad => N_58169,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_25_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(82),
cin => N_57464);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_25_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57466,
datad => N_58146,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_26_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(83),
cin => N_57468);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_26_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57470,
datad => N_58123,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_27_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(84),
cin => N_57472);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_27_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57474,
datad => N_58100,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_28_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(85),
cin => N_57476);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_28_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57478,
datad => N_58077,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_29_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(86),
cin => N_57480);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_29_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57482,
datad => N_58054,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_30_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(87),
cin => N_57484);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_30_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57486,
datad => N_58031,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_31_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(88),
cin => N_57488);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_31_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57490,
datad => N_58008,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_32_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(89),
cin => N_57492);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_32_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57494,
datad => N_57985,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_33_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(90),
cin => N_57496);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_33_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57498,
datad => N_57962,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_34_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(91),
cin => N_57500);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_34_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57502,
datad => N_57939,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_35_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(92),
cin => N_57504);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_35_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57506,
datad => N_57916,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_36_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(93),
cin => N_57508);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_36_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57510,
datad => N_57893,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_8_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(65),
cin => N_57512);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_8_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57514,
datad => N_57870,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_9_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(66),
cin => N_57516);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_9_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57518,
datad => N_57847,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_10_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(67),
cin => N_57520);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_10_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57522,
datad => N_57824,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_11_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(68),
cin => N_57524);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_11_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57526,
datad => N_57801,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_12_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(69),
cin => N_57528);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_12_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57530,
datad => N_57778,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_13_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(70),
cin => N_57532);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_13_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57534,
datad => N_57755,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_14_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(71),
cin => N_57536);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_14_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57538,
datad => N_57732,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_15_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(72),
cin => N_57540);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_15_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57542,
datad => N_57709,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_16_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(73),
cin => N_57544);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_16_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57546,
datad => N_57686,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_17_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(74),
cin => N_57548);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_17_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57550,
datad => N_57663,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_18_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(75),
cin => N_57552);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_18_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57554,
datad => N_57640,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_19_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(76),
cin => N_57556);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_19_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57558,
datad => N_57617,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_20_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(77),
cin => N_57560);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_20_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57562,
datad => N_57594,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_21_Z_CARRY_3_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(78),
cin => N_57564);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_21_Z_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_57566,
datad => N_57571,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_2_IV_0_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"0ee0eeee0ee0eaea")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_IV_0\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4233\,
datae => \GRLFPC2_0.FPI.LDOP\,
datad => \GRLFPC2_0.FPI.OP2\(63),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(22),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4534\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(12),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIHTQC5_20_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"f0f05041f0f05050")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(20),
datae => \GRLFPC2_0.FPI.LDOP_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6_I\,
datac => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_10: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"faf5f9f9af5f9f9f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_10\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10879\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10865\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10866\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(1),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10878\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_236_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"0f00c4c40f008080")
port map (
combout => N_36149,
dataf => \GRLFPC2_0.FPO.EXP\(8),
datae => \GRLFPC2_0.FPI.LDOP\,
datad => \GRLFPC2_0.FPI.OP2\(60),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(249),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_45_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"ffffa0a03000a0a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2779\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83),
datad => N_32048_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2671\,
datab => N_33043_I,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85),
datag => N_33001_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_234_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"0f00c4c40f008080")
port map (
combout => N_36203,
dataf => \GRLFPC2_0.FPO.EXP\(10),
datae => \GRLFPC2_0.FPI.LDOP\,
datad => \GRLFPC2_0.FPI.OP2\(62),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(247),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_235_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"0f00c4c40f008080")
port map (
combout => N_36176,
dataf => \GRLFPC2_0.FPO.EXP\(9),
datae => \GRLFPC2_0.FPI.LDOP\,
datad => \GRLFPC2_0.FPI.OP2\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(248),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"f00ff00f88778877")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(226),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"f00ff00f88778877")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(227),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"f00ff00f88778877")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(229),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"f00ff00f88778877")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(225),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_9_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"ffccffdcffecffdc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_10\,
dataf => N_31999_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85),
datad => N_32210,
datac => N_32206_2,
datab => N_32712_3,
dataa => N_31767_2,
datag => N_32705_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_22_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"9a95a5a59a955555")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(22),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(209),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"f00ff00f88778877")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(228),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"9a95a5a59a955555")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(19),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(212),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(55),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(176),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_X2_RNIKKUG2_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"0f00808000008080")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
datae => N_32908_1,
datad => N_33136_1,
datac => N_32487_2,
datab => N_28591_1,
dataa => N_28580_1,
datag => N_32394_I);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_41_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(41),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(190),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"00f0080800f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_6\,
dataf => N_32131_1,
datae => N_31819_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datab => N_32136_2,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(78),
datag => N_32567_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(8),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(223),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_6_1_RNIHVHV_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"c0000a0ac0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_0_0\,
dataf => N_31838_1,
datae => N_31766_1,
datad => N_27553_1,
datac => N_31788,
datab => N_32775_1,
dataa => N_31725_1,
datag => N_33176);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(28),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(203),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(50),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(181),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_20_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(20),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(211),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_9_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(9),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(222),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_44_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(44),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(187),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_12_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(12),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(219),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"f6f9f9f96f9f9f9f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10889\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10869\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5343\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10882\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_0_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"0ffff7f7fffff7f7")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_0\(47),
dataf => N_32142_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(78),
datab => N_27929_1,
dataa => N_31865_1,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"000a808000008080")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datae => N_31996_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(81),
datac => N_31808_1,
datab => N_27553_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(78),
datag => N_32662_I);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_49_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(49),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(182),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_GEN: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"0f00ec800000ec80")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.GEN\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10579\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(372),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(371),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(314),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(114));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_24_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(24),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(207),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_3_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"0555fdfd0fffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_3\(47),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
datae => N_31715_1,
datad => N_31769_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(78),
dataa => N_31999_1,
datag => N_32142_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(51),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(180),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_46_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(46),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(185),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_11_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"f0004c4cf0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_2\,
dataf => N_33138_1,
datae => N_31775_1,
datad => N_31766_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85),
datab => N_31765_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83),
datag => N_31763_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(178),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_43_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(43),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(188),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(33),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(198),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"c000a0a0c0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_2\,
dataf => N_32627_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
datad => N_33136_2,
datac => N_32069_2,
datab => N_31996_1,
dataa => N_28580_1,
datag => N_32032_I);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"50001000a0a02020")
port map (
combout => N_52474,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82),
datac => N_32220_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(81),
datag => N_32567_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_38_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(38),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(193),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(31),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(200),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(25),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(206),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(48),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(183),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_42_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(42),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(189),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"f0000808f0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_0\,
dataf => N_32069_2,
datae => N_31919_1,
datad => N_33057_1,
datac => N_31768_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
datag => N_31718_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_14_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(14),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(217),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(32),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(199),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_30_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(30),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(201),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_10_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(10),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(221),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_45_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(45),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(186),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_35_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(35),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(196),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(52),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(179),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_39_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(39),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(192),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_9_0_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"f0ffffff70775757")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_9_0\(31),
dataf => N_32739,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datad => N_32705_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84),
datab => N_31940_1,
dataa => N_32487_2,
datag => N_33298);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(54),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(177),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(47),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(184),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(17),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(214),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(224),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(18),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(213),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(26),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(205),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(13),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(218),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(34),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(197),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_15_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(15),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(216),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_23_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(23),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(208),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(11),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(220),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_40_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(40),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(191),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(27),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(204),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(56),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(175),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_17_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"0000b3ff70f077ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_17\(47),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83),
datae => N_32619_1,
datad => N_31715_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
datab => N_32128_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84),
datag => N_28580_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(36),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(195),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(29),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(202),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_21_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(21),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(210),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"0000202000f02020")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_4\,
dataf => N_32885_I,
datae => N_31763_1,
datad => N_33138_1,
datac => N_32708_2,
datab => N_32688_1,
dataa => N_31767_2,
datag => N_31775_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"1010404010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_2\,
dataf => N_31765_1,
datae => N_32066_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85),
datac => N_31839_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_37_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(37),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(194),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_16_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(16),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(215),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"ccccccccfccccdcd")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_11\,
dataf => N_32739,
datae => N_33298,
datad => N_32632_1,
datac => N_32673_I,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85),
datag => N_32050_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_9_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"00f0080000000800")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_3\,
dataf => N_31769_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(78),
datab => N_31808_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(81),
datag => N_31941_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_I_1_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"5f5f7fffffff7fff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_1\(31),
dataf => N_31941_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79),
datac => N_32775_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\(78),
datag => N_32070_1);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN17_SHDVAR: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"0000000000050101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN17_SHDVAR\,
dataf => N_59196,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
dataa => N_59195,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a80aa0a008080000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_1\,
dataf => N_32120_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datac => N_31921_1,
datab => N_33314_4,
dataa => N_31924_1,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_8_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"1000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2639\,
dataf => N_31762_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84),
datac => N_32032_I,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\(78),
datag => N_31921_1_0);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_1_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"0080a0a000000000")
port map (
combout => N_32196,
dataf => N_31723_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(81),
datac => N_31999_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83),
dataa => N_32705_1,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A20_1_RNIRNDAC_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"00000000f0006000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datad => N_31766_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datag => N_32140_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_13_C_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"cfcfffccefefffec")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_13_C\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(74),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(76),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_377\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(63),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(71));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_120_RNI3H4S: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"fefafefabafabafa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10927_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(49),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_27_S_0_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10918_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0\,
datag => N_55054_RETO);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CARRY_0_BUF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ff00")
port map (
cout => N_81973,
datad => VCC,
cin => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff2000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_13\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_7\,
datae => N_32841,
datad => N_32141_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A28_24_0\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_1_RNIDHHS: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"d0ddfdff2f220200")
port map (
combout => N_34177,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10634\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10635\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(316));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00000080")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_1\,
dataf => N_32994,
datae => N_32052_1,
datad => N_32688_1,
datac => N_31769_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_20_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0c0cfc0c0c0c0c")
port map (
combout => N_80614,
dataf => N_81711,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_7__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_8__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_9\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_20_RNO_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000ff0ff")
port map (
combout => N_81711,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_14__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10070\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10130\,
datac => N_76344);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_11_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"2222222e22222222")
port map (
combout => N_80619,
dataf => N_81709,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_11__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_15__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_17__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_10\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_11_RNO_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ffff00ffff")
port map (
combout => N_81709,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10077\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10137\,
datad => N_76344);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_127_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"707f0000f0ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2462\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV\,
datae => N_81707,
datad => N_79923,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN10_FEEDBACK\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(48));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_127_RNO_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000f00000")
port map (
combout => N_81707,
dataf => N_79937,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748\,
datac => N_56);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_1_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751_RETI\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G0_I_0_2_RETI\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G0_I_0_RETI\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0707070505070505")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
dataf => N_26592,
datae => N_26591,
datad => N_26534,
datac => N_81690,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_I\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA_SUB: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff3fffffffffff")
port map (
combout => N_81690,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
datae => \GRLFPC2_0.FPI.LDOP_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN1_CCIN_RNI5VI831: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fef1fff1fefeffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN25_NOTPROP\,
datae => N_81684,
datad => N_81301,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SBLSBS_1\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_959_I\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_10_RNIIGE42_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ccccf000cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(11),
dataf => N_81674,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_20\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_10\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_12_RNI8U5B_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fffffffffffffff")
port map (
combout => N_81674,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_13\(11),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_12\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_2\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_3\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNILSA9U_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffccf0ccffccffcc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(13),
dataf => N_81640,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_8\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_7\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O17_4_RNIHBO7L_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000f00ff")
port map (
combout => N_81640,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_12\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A17_0\(13),
datad => N_33206,
datac => N_33193);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNI7IDRJ_12_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00f0f0fffff0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(12),
dataf => N_81634,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_9_RNIATI07_12_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000f")
port map (
combout => N_81634,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_7\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2311\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_RNO_10_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"55dd77ff50d872fa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(10),
dataf => N_81630,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(10),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_RNO_0_10_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000f0ff0fffff")
port map (
combout => N_81630,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(10),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_11_RNIFI642: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffeaaaffffaaa8")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5330\,
dataf => N_81626,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\(11),
datad => \GRLFPC2_0.FPO.EXP\(10),
datac => \GRLFPC2_0.FPO.EXP\(9),
datab => \GRLFPC2_0.FPO.EXP\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_RNO_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff0cfff3ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(46),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(11),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A28_31_1_RNI6JCVK_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffff00ff20")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_12\,
dataf => N_81621,
datae => N_28591_1,
datad => N_33201,
datac => N_31766_1,
datab => N_31996_1,
dataa => N_32418_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_12_RNIJ8PGA_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffff0ffffff00")
port map (
combout => N_81621,
dataf => N_33207_1,
datae => N_33208,
datad => N_33196,
datac => N_32221_1);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_5_RNI6DKJ: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ffffffffffffff")
port map (
combout => N_81619,
dataf => \GRLFPC2_0.FPO.EXP\(7),
datae => \GRLFPC2_0.FPO.EXP\(6),
datad => \GRLFPC2_0.FPO.EXP\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_RNO_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"efabcd8967234501")
port map (
combout => N_59307,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(2),
datac => N_81615,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_RNO_0_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00ff00ff")
port map (
combout => N_81615,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datae => N_59228,
datad => N_59226);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNISLF71_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"45badf20ba4520df")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_58\(56),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_1\,
datad => N_81611,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10634\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10635\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_0_RNI1K3E_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f0ff0fffffffff")
port map (
combout => N_81611,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5771\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000fffc3f3c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(11),
dataf => N_81609,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_SUB_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"001040500a1a4a5a")
port map (
combout => N_81609,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(9),
datae => N_59191,
datad => N_59217,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_RNITJ5N_40_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"5555ccccff00f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(15),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => N_59263,
datac => N_59262,
datab => N_59246,
dataa => N_81599);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNI6PS3_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff00ff0000ffff")
port map (
combout => N_81599,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_RNISF5N_40_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0ff005555cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(17),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => N_59263,
datac => N_59272,
datab => N_59246,
dataa => N_81599);
GRLFPC2_0_FPI_LDOP: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0000")
port map (
combout => \GRLFPC2_0.FPI.LDOP\,
dataf => \GRLFPC2_0.R.MK.RST\,
datae => N_81563);
GRLFPC2_0_FPI_LDOP_SUB: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffdfff55ff55ff55")
port map (
combout => N_81563,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7612_I_A7_10\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7612_I_A7_6\,
datad => \GRLFPC2_0.R.MK.RST2\,
datac => \GRLFPC2_0.R.STATE_O_3\(0),
datab => \GRLFPC2_0.R.STATE_O_3\(1),
dataa => N_7);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIB1PT_10_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ffaaaaccccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(14),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datad => N_81561,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNI9QTC_244_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff00ff0000ffff")
port map (
combout => N_81561,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_RNO_12_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00fff0f0aaaacccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(12),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datad => N_81559,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_RNO_0_12_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff00ff0000ffff")
port map (
combout => N_81559,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN26_NOTAINFNAN: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff800000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7144\,
dataf => N_81507,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN26_NOTAINFNAN_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN26_NOTAINFNAN_SUB: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fffffffffffffff")
port map (
combout => N_81507,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(243),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(237));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0cccc0f00cccc")
port map (
combout => N_80625,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10076\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10136\,
datac => N_76344,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_2_RNO_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000001b")
port map (
combout => N_81263,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_10__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_13__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_16__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10080\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10140\,
dataa => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIBKAH_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0cccc0f00cccc")
port map (
combout => N_80635,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10027\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10087\,
datac => N_76344,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0cccc0f00cccc")
port map (
combout => N_80674,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10082\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10142\,
datac => N_76344,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_141_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0aff0a00caffca00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(141),
dataf => N_59283,
datae => \GRLFPC2_0.FPO.FRAC\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
datac => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(143));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_7_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000020000000000")
port map (
combout => N_33203,
dataf => N_31996_1,
datae => N_32064_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_13_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000100000000000")
port map (
combout => N_33209,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(81),
datae => N_33176,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_12_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030303010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2306\,
dataf => N_33314_4,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(81),
datad => N_31715_1,
datac => N_31924_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_48_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"4000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2042\,
dataf => N_32131_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(81),
datad => N_31762_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_5_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff005f00ff007f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_5\(11),
dataf => N_31766_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(81),
datad => N_32064,
datac => N_32047_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_RNIFLE5A_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0040000000510000")
port map (
combout => N_33196,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(81),
datae => N_31769_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN13_GEN: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"2d002000d2000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN13_GEN\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SALSBS_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5446\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(370));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_12_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000040")
port map (
combout => N_33208,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(81),
datae => N_33176,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_A26_17_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0400000000000000")
port map (
combout => N_32064,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3363c3633c6ccc6c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10944\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(241));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_RNI20S01_68_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0ccfff0f0cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(68),
datae => \GRLFPC2_0.FPI.LDOP_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(68),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(68));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3ccccccc6c6c6c6c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(239));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_122_RNIJ6N64_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f0f0f0ff0f0f0f")
port map (
combout => N_81301,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SCLSBS_2\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0f0f03030f0303")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897\,
dataf => N_26592,
datae => N_26591,
datad => N_26534,
datac => N_81293,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_SUB: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff03ffff0303ffff")
port map (
combout => N_81293,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_0_RNO_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000001b")
port map (
combout => N_81259,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_7__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_4__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_3__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10074\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10134\,
dataa => N_76344);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_2_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcfcfc0cfcfcfcfc")
port map (
combout => N_80624,
dataf => N_81263,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_4__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_6__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
datab => N_79982);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_0_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0c0cfc0c0c0c0c")
port map (
combout => N_80631,
dataf => N_81259,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_6__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_5__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7782_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNI032Q_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0cccc0f00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10081\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10141\,
datac => N_76344,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333331131313131")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10026\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.NOTPROP_3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN25_GEN\,
datac => N_59288,
datab => N_81250,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_SUB_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f00ff000ff0fff")
port map (
combout => N_81250,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0c0c04040c0404")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
dataf => N_26592,
datae => N_26591,
datad => N_26534,
datac => N_81248,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_SUB: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000100010001")
port map (
combout => N_81248,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\,
datad => \GRLFPC2_0.FPI.LDOP_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNI93GF6U1_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfcfc0c0cfc0cfc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(1),
dataf => N_26534,
datae => N_26586,
datad => N_26585,
datac => N_81224,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNI47VJL01_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30303f3f303f303f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(0),
dataf => N_26534,
datae => N_26588,
datad => N_26587,
datac => N_81224,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNINUA3_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000ff0000")
port map (
combout => N_81224,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIEH8TUC2_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfcfc0c0cfc0cfc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(2),
dataf => N_26534,
datae => N_26584,
datad => N_26583,
datac => N_81224,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIJO44BK2_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfcfc0c0cfc0cfc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(3),
dataf => N_26534,
datae => N_26582,
datad => N_26581,
datac => N_81224,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_3_1_RNI1994A_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"8000000000000000")
port map (
combout => N_32497,
dataf => N_32070_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_13_1_RNIQDR1A_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0048000000000000")
port map (
combout => N_33201,
dataf => N_31996_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_8_RNO_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000020002020")
port map (
combout => N_32046,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(81),
datae => N_31788,
datad => N_32022_I,
datac => N_31989_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_9_RNO_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0003000a000200")
port map (
combout => N_32048,
dataf => N_31724_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(81),
datad => N_32048_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_RNIPC1Q1_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f232202020202020")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_2_1_CO1\,
dataf => N_81177,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10634\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(316));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIV4B41_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff000ff0ff0ff00")
port map (
combout => N_81177,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN_RNIFOI51_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00aaaa0f0fcccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(9),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\(5),
datac => N_81171,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNI7QTC_243_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff00ff0000ffff")
port map (
combout => N_81171,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(243));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIRKAF2_16_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffc000c0ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(31),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIS5NO1_247_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff800000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1919\,
dataf => N_81152,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_I_0_A2_4\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(247),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(248),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(249));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIJ28I_250_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fffffffffffffff")
port map (
combout => N_81152,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(251),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(253),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(250),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(257));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_59_RNIS8B41: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00f0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO_0\,
datae => \GRLFPC2_0.FPI.LDOP_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(100),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(100),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(100));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_19_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"4000500040000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5394_RETI\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(58),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_317__G1\,
dataa => \GRLFPC2_0.FPI.LDOP_4\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIE0BH_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0cccc0f00cccc")
port map (
combout => N_80634,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10026\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10086\,
datac => N_76344,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_RNIQKGK41_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"98ff980010ff1000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_57__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10085\,
datad => N_76344,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"4c4c4c44444c4444")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4534\,
dataf => N_26592,
datae => N_26591,
datad => N_26534,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_I\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_A26_9_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"4800000000000000")
port map (
combout => N_32056,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(81),
datae => N_31723_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_43_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ff0000f0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(43),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(72),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datad => \GRLFPC2_0.FPI.LDOP_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(72));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN5_ZERO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"77770fffeeeefff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffa0ff8000a00080")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(18),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffa0ff8000a00080")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(17),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_30_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffa000a0ff800080")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(30),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffa000a0ff800080")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(29),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_RNI94S01_76_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0ccfff0f0cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(76),
datae => \GRLFPC2_0.FPI.LDOP_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(76),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(76));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_RNI94S01_74_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0ccfff0f0cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(74),
datae => \GRLFPC2_0.FPI.LDOP_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(74),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(74));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_RNIHH821_98_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0fff0ccf000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(98),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO_0\,
datad => \GRLFPC2_0.FPI.LDOP_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(98),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(98));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_RNI20S01_95_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0fff0ccf000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(95),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO_0\,
datad => \GRLFPC2_0.FPI.LDOP_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(95),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(95));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_RNIH0S01_97_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0fff0ccf000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(97),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO_0\,
datad => \GRLFPC2_0.FPI.LDOP_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(97),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(97));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_RNI00S01_94_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0fff0ccf000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(94),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO_0\,
datad => \GRLFPC2_0.FPI.LDOP_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(94),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(94));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaacc00aaaac000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaacc00aaaac000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(8),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaacc00aaaac000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_12_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffa000a0ff800080")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(12),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaacc00aaaac000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffa000a0ff800080")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(11),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_10_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffa000a0ff800080")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(10),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_9_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffa000a0ff800080")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(9),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_16_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffa0ff8000a00080")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(16),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaacc00aaaac000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_15_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffa000a0ff800080")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(15),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaacc00aaaac000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaacc00aaaac000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(13),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_14_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffa000a0ff800080")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(14),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_76_RNIRGB41: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ccccff00f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO_0\,
datae => \GRLFPC2_0.FPI.LDOP_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(101),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(101),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(101));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_86_RNI7HB41: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ccccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
dataf => \GRLFPC2_0.FPI.LDOP_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(105),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(105),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(105));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_108_RNIOUO51: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ccccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
dataf => \GRLFPC2_0.FPI.LDOP_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(86),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(86),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(86));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_84_RNI5TB41: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ccccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
dataf => \GRLFPC2_0.FPI.LDOP_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(80));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_95_RNIROB41: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ccccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
dataf => \GRLFPC2_0.FPI.LDOP_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(106),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(106),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(106));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_120_RNIC6P51: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ccccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
dataf => \GRLFPC2_0.FPI.LDOP_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(84));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_92_RNIU4C41: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ccccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
dataf => \GRLFPC2_0.FPI.LDOP_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(81));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_78_RNI0LB41: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ccccff00f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO_0\,
datae => \GRLFPC2_0.FPI.LDOP_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(103),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(103),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(103));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_117_RNIL6P51: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ccccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
dataf => \GRLFPC2_0.FPI.LDOP_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(85));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_80_RNIRGB41: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ccccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
dataf => \GRLFPC2_0.FPI.LDOP_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(104),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(104),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(104));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_9_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_9__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10073\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10133\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_18__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10064\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10124\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIR0CD_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_19__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10063\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10123\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_20_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_20__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10062\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10122\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNID0AD_21_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_21__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10061\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10121\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIF8AD_22_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_22__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10060\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10120\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIHGAD_23_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_23__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10059\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10119\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIJOAD_24_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_24__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10058\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10118\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIL0BD_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_25__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10057\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10117\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_26__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10056\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10116\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_27__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10055\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10115\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_28__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10054\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10114\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_29__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10053\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10113\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_30_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_30__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10052\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10112\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_31__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10051\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10111\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_32__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10050\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10110\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_33__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10049\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10109\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_34__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10048\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10108\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_35_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_35__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10047\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10107\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_36__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10046\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10106\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_37_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_37__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10045\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10105\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_38_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_38__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10044\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10104\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_39_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_39__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10043\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10103\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_40_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_40__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10042\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10102\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_41_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_41__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10041\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10101\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_42_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_42__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10040\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10100\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_43_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_43__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10039\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10099\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_44_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_44__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10038\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10098\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_45_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_45__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10037\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10097\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_46_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_46__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10036\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10096\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_47__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10035\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10095\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_48__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10034\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10094\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_49_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_49__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10033\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10093\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_50__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10032\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10092\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIJ0AD_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_51__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10031\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10091\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_52__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10030\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10090\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNINGAD_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_53__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10029\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10089\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIPOAD_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_54__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10028\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10088\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_9_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80673,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_9__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80672,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_18__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNI7LTG_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80671,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_19__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_20_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80670,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_20__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_3_RNIIKQG: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80669,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_21__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIM0RG_22_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80668,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_22__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIPCRG_23_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80667,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_23__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNISORG_24_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80666,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_24__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIV4SG_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80665,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_25__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80664,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_26__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80663,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_27__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80662,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_28__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_80661,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_29__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_30_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_80660,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_30__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_80659,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_31__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_80658,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_32__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_80657,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_33__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80656,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_34__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_35_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80655,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_35__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80654,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_36__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_37_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80653,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_37__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_38_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80652,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_38__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_39_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80651,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_39__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_40_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80650,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_40__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_41_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80649,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_41__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_42_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80648,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_42__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_43_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80647,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_43__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_44_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80646,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_44__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_45_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80645,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_45__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_46_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80644,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_46__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_80643,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_47__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_80642,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_48__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_49_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_80641,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_49__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_80640,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_50__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIV39H_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_80639,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_51__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_80638,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_52__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_RNI5S9H: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_80637,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_53__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNI88AH_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_80636,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_54__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNICGGO41_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80633,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_57__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80632,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_3__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_10_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80630,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_10__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_16_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80629,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_16__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80627,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_13__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80626,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_4__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_15_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80623,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_15__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80622,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_5__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80621,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_11__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80620,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_17__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80618,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_7__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80617,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_8__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_14_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_80615,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_14__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_101_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaff00f0f0cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(101),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datad => \GRLFPC2_0.FPO.FRAC\(14),
datac => \GRLFPC2_0.FPO.FRAC\(12),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_100_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaff00f0f0cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(100),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datad => \GRLFPC2_0.FPO.FRAC\(15),
datac => \GRLFPC2_0.FPO.FRAC\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_77_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaff00f0f0cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(77),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(38),
datac => \GRLFPC2_0.FPO.FRAC\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_99_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaff00f0f0cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(99),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datad => \GRLFPC2_0.FPO.FRAC\(16),
datac => \GRLFPC2_0.FPO.FRAC\(14),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A3_5_SUB_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff00")
port map (
combout => N_79998_RETO,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2462_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_4_0_RETO\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(73));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_98_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(98),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_RETO\,
datad => \GRLFPC2_0.FPO.FRAC_RETO\(17),
datac => \GRLFPC2_0.FPO.FRAC_RETO\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(98),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(40));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_97_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(97),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_RETO\,
datad => \GRLFPC2_0.FPO.FRAC_RETO\(18),
datac => \GRLFPC2_0.FPO.FRAC_RETO\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(97),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_76_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(76),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_RETO\,
datad => \GRLFPC2_0.FPO.FRAC_RETO\(39),
datac => \GRLFPC2_0.FPO.FRAC_RETO\(37),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(76),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_95_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(95),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_RETO\,
datad => \GRLFPC2_0.FPO.FRAC_RETO\(20),
datac => \GRLFPC2_0.FPO.FRAC_RETO\(18),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(95),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_74_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaff00f0f0cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(74),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_RETO\,
datad => \GRLFPC2_0.FPO.FRAC_RETO\(39),
datac => \GRLFPC2_0.FPO.FRAC_RETO\(41),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(74),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_94_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(94),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_RETO\,
datad => \GRLFPC2_0.FPO.FRAC_RETO\(21),
datac => \GRLFPC2_0.FPO.FRAC_RETO\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(94),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_92_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(92),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_RETO\,
datad => \GRLFPC2_0.FPO.FRAC_RETO\(23),
datac => \GRLFPC2_0.FPO.FRAC_RETO\(21),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(92),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_91_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(91),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_RETO\,
datad => \GRLFPC2_0.FPO.FRAC_RETO\(24),
datac => \GRLFPC2_0.FPO.FRAC_RETO\(22),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(91),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_68_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(68),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_RETO\,
datad => \GRLFPC2_0.FPO.FRAC_RETO\(47),
datac => \GRLFPC2_0.FPO.FRAC_RETO\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(68),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_90_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(90),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_RETO\,
datad => \GRLFPC2_0.FPO.FRAC_RETO\(25),
datac => \GRLFPC2_0.FPO.FRAC_RETO\(23),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(90),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_89_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(89),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_RETO\,
datad => \GRLFPC2_0.FPO.FRAC_RETO\(26),
datac => \GRLFPC2_0.FPO.FRAC_RETO\(24),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(89),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_88_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(88),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_RETO\,
datad => \GRLFPC2_0.FPO.FRAC_RETO\(27),
datac => \GRLFPC2_0.FPO.FRAC_RETO\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(88),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_87_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(87),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_RETO\,
datad => \GRLFPC2_0.FPO.FRAC_RETO\(28),
datac => \GRLFPC2_0.FPO.FRAC_RETO\(26),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(87),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccff00f0f0aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(60),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_RETO\,
datad => \GRLFPC2_0.FPO.FRAC_RETO\(53),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_176__G2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(60));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccff00f0f0aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(59),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_RETO\,
datad => \GRLFPC2_0.FPO.FRAC_RETO\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_175__G2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(59));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_72_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0ccffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0_RETO\(72),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(72),
datad => N_26534_RETO,
datac => N_26564_RETO,
datab => N_26563_RETO);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_72_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000f0ccf0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1_RETO\(72),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(14),
datad => N_26534_RETO,
datac => N_26560_RETO,
datab => N_26559_RETO);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_5_2_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"88ff888888ff88f8")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_5_1_RETO\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2466_1_RETO\,
dataa => N_28949_RETO);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_12_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0033003300330f33")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_455_RETO\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(4),
datab => N_28949_RETO);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A3_10_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2463_RETO\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_13_1_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00c000c000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_1\,
datad => CPI_D_INST_RETO(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_377_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_13_C_RETO\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_1_RNI1GKU1_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000dd000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_I_0_0_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_RETO\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5330_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_26_RNI5C422_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000fa0033")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_I_0_0_RETO\,
datac => \GRLFPC2_0.FPO.FRAC_RETO\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0_RETO\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A2_2_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"2200222222002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_2_RETO\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2474_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1164_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_88_RNIEU7R: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff3")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(77),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_237_RETO\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_231_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(231),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(231));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_15_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(15),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_15__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(15));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_13_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"1113113313133333")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G1_1_RETI\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(374),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(12),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(231));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_22_RNIGNLN: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_RETO\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_79_RNIKRLN: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO\(55),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_38_RNIFRLN_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO\(54),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A3_5_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffffffdf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO\,
dataf => N_79998_RETO,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_78_RNIJRLN: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_77_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(77),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(77),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(77));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_99_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(99),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(99),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(99));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_89_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(89),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(89),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(89));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_88_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(88),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(88),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(88));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_92_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(92),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(92),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(92));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_RNI6S5J_77_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(77),
datae => \GRLFPC2_0.FPI.LDOP_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(77));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_91_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(91),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(91),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(91));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_90_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(90),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(90),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(90));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_RNI7O5J_99_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(99),
datae => \GRLFPC2_0.FPI.LDOP_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(99));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_87_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(87),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(87),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(87));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_RNI106J_88_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(88),
datae => \GRLFPC2_0.FPI.LDOP_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(88));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_RNI906J_89_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(89),
datae => \GRLFPC2_0.FPI.LDOP_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(89));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_RNIRN5J_92_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(92),
datae => \GRLFPC2_0.FPI.LDOP_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(92));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_RNION5J_91_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(91),
datae => \GRLFPC2_0.FPI.LDOP_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(91));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_RNIQ36J_90_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(90),
datae => \GRLFPC2_0.FPI.LDOP_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(90));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_RNI106J_87_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(87),
datae => \GRLFPC2_0.FPI.LDOP_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(87));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIHOAD_14_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_14__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10068\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10128\,
datad => N_76344);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_5_RNI1VPN: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f0f0ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
dataf => \GRLFPC2_0.FPI.LDOP_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(113),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_372__G1_RETO\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_RNIK2NQ_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0ff0000f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(59),
datae => \GRLFPC2_0.FPI.LDOP_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_318__G1_RETO\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0fffffff000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(60),
datae => \GRLFPC2_0.FPI.LDOP_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_319__G1_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_21_RNIM4491: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000aaf00000aacc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(114),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_RETO\,
datae => \GRLFPC2_0.FPI.LDOP_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1_RETO\(114),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0_RETO\(114),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_3_I_RETO\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_115_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000f0000000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(115),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_RETO\,
datae => \GRLFPC2_0.FPI.LDOP_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1_RETO\(115),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0_RETO\(115));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_12_RNIK9SJ1_8: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000fffc0200fefc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(65),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIB0AD_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_11__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10071\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10131\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNINGBD_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_17__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10065\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10125\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIJ0BD_15_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_15__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10067\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10127\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_72_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfcfcfc0c0cfc0c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(72),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1_RETO\(72),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0_RETO\(72),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(72));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_4_RNIFUIF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(72),
datae => \GRLFPC2_0.FPI.LDOP_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(72));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_BUSYMULXFF_UN2_TEMP: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"dddfdddddddfdddf")
port map (
combout => \GRLFPC2_0.FPO.BUSY_O\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3924_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.BUSYMULXFF.UN2_TEMP_2_RETO\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"1111555555055555")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_217_RETO\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(4),
datab => CPI_D_INST_RETO(6),
dataa => N_79941_RETO);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIL8BD_16_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_16__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10066\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10126\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIFGAD_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_13__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10069\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10129\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNI9O9D_10_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_10__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10072\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10132\,
datad => N_76344);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RET_0_RNI045R: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"08f80808f4040404")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_I_I_0_RETO\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.U_RDN_1_RETO\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.UN17_U_RDN_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.TEMP_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_RETO\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_RETO\(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RET_1_RNI2H931: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I_RETO\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_5_3_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffa0808080")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_5_2_RETO\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_5_1_RETO\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_0\,
datac => CPI_D_INST_RETO(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_377_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_13_C_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A2_3_2_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3cccffff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_2_RETO\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2466_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(81));
GRLFPC2_0_COMB_V_MK_BUSY_2_4_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.FPO.BUSY_O_0\,
dataf => \GRLFPC2_0.FPO.BUSY_O\,
datae => RST_RETO);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_5_1_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000220255557757")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2809_1_RETO\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_217_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_0\,
datad => CPI_D_INST_RETO(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_377_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2457_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(73));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_12_RNIJ9FU_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf0fcfcfefafefe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0_4__G0_2_RETO\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_217_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_455_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2555_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_4_0_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A2_3_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"4040404040404000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2463_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2462_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_4_0_RETO\(4),
datac => N_31763_1_RETO,
datab => N_31723_1_RETO,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_255_RETO\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNILTUK_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_7__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10135\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIFTUK_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_4__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10078\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10138\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIJTUK_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_6__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10076\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10136\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIHTUK_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_5__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10077\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10137\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIDTUK_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_3__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10079\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10139\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNINTUK_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_8__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10074\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10134\,
datad => N_76344);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(8),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_8__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(8));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNIMA9E3_14_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0103050f113355ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349_I_0_RETI\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_DIVMULTV\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(14));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_43_RNI3VGR1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0033003000220020")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO\(53),
datac => N_28952_RETO,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO\(84),
dataa => CPI_D_INST_RETO(12));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_40_RNISUGR1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0033003000220020")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO\(54),
datac => N_28951_RETO,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO\(6),
dataa => CPI_D_INST_RETO(8));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_35_RNI7VGR1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0033003000220020")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO\(55),
datac => N_28950_RETO,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO\(79),
dataa => CPI_D_INST_RETO(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_31_RNI8JF23: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f0c0a08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO\,
datab => N_28945_RETO,
dataa => CPI_D_INST_RETO(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_27_RNIRFV53: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f0c0a08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO\(2),
datab => N_28947_RETO,
dataa => CPI_D_INST_RETO(7));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_23_RNI3DNN2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff003caabe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(82),
dataa => CPI_D_INST_RETO(11));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_15_RNITQGR1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0033003000220020")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO\(1),
datac => N_28946_RETO,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_RETO\,
dataa => CPI_D_INST_RETO(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_5_1_RNIIU4N_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf0fcf0fcf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0_4__G0_4_RETO\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2809_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_5_2_RETO\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_729_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_13_1_RNIHC652_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff10")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0_4__G0_4_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0_4__G0_2_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNIHRCES_9_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f00ff0f0fffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G0_I_0_RETI\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(374),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_14_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(14),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_14__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(14));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_1_RNO_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"01330133013305ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G0_I_0_2_RETI\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(375),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_DIVMULTV\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(14));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_9_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(9),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_16_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(10),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_16__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"faaaf000feeefccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_RETI\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(375),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_142_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(142),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_14\(142),
datae => \GRLFPC2_0.FPO.FRAC\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_RNI8CIC: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00000000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G0_I_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349_I_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIKLTU_230_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000377700003fff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G0_0_O2_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(374),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5394\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(12),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(230),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_18_RNI8A8I1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"dc50ffff23af0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5391\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G0_0_O2_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349_I_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_13_RNI8RTQ: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff737773008c888c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5410\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G1_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349_I_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN2_NOTDECODEDUNIMP_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000050105050")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.STARTSHFT.UN2_NOTDECODEDUNIMP_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1902\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19\(45),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(66),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(67),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(64));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00600000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_0\,
datae => N_32340_1,
datad => N_33298,
datac => N_32786_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_10_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000feff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_10\(11),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_0\(11),
datae => N_32049,
datad => N_33071_1,
datac => N_33232,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_4_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f7ffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_4\(47),
dataf => N_32628,
datae => N_32645_3,
datad => N_32124_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
datab => N_32645_2,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff9000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_17\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_10\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_0_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(81),
datac => N_32243,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_49_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0200")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_6\,
dataf => N_32350,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_31_1\(48),
datac => N_31989_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A3_RNIB5IE9_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff000040c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_0\,
datae => N_32340_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2546\,
datab => N_31819_2,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff4000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_16\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_1\,
datae => N_32199,
datad => N_32708_2,
datac => N_32221_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_45_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff909090ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2_0\,
dataf => N_33138_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2513\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2499\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2538\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_10_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f8f0f0f088000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_4\,
dataf => N_32413_2,
datae => N_32400,
datad => N_32272_2,
datac => N_31838_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_A30_12_1_RNISUNR4_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffff00ff10")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2_2\,
dataf => N_33148,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_255\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2784\,
datac => N_31931_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
GRLFPC2_0_COMB_UN2_HOLDN_0_A3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"4000000000000000")
port map (
combout => \GRLFPC2_0.N_1470\,
dataf => \GRLFPC2_0.COMB.UN2_HOLDN_0_A3_13\,
datae => \GRLFPC2_0.COMB.UN2_HOLDN_0_A3_11\,
datad => \GRLFPC2_0.COMB.UN2_HOLDN_0_A3_10\,
datac => \GRLFPC2_0.COMB.V.E.FPOP_1\,
datab => \GRLFPC2_0.FPCI_O\(62),
dataa => \GRLFPC2_0.FPCI_O\(69));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_2_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0bffffffbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_2\(11),
dataf => N_32032_I,
datae => N_33057_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(81),
datac => N_31715_1,
datab => N_31718_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_0_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ddddddd0fffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_0\(11),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_A26_6_1\(11),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_A26_23_0\(11),
datad => N_32070_1,
datac => N_31864_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_63_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff444fffff000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_346\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1810\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_9_0\(62),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2490\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_63_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0b00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1812\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2494\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_247\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0080")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_12\,
dataf => N_33067,
datae => N_33060,
datad => N_32124_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(81),
datab => N_32485_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff1000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_7\,
dataf => N_32785,
datae => N_32273,
datad => N_31996_1,
datac => N_32220_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff10")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_16\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_8\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_7\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_6\,
datac => N_33145_4,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_10_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff10")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_8\,
dataf => N_32699,
datae => N_32708,
datad => N_32698,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_1_1\(58),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff8000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_15\,
dataf => N_32693,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_8\,
datad => N_32290_1,
datac => N_32673_I,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0b0b0bff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_6\,
dataf => N_32198_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_12_0\(57),
datad => N_32207_1,
datac => N_32232,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff4000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_13\,
dataf => N_32427,
datae => N_32432,
datad => N_32413_2,
datac => N_32394_I,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff1f110f00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_9\,
dataf => N_32768,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A24_8_1\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A24_10_1\(55),
datac => N_33298,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff1000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_10\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_0\,
datae => N_32558,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_44_0\(54),
datac => N_32220_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_49_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff8000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_13\,
dataf => N_32348,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_4\,
datad => N_32344_1,
datac => N_32327,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_41_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffff111f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_41__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1788\,
datae => N_33271,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2689\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2526\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_1_0_39_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff909090ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_1_0\(39),
dataf => N_31925_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2666\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2538\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2652\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_9\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_0\,
datae => N_31993,
datad => N_31983,
datac => N_33040,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff10")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_7\,
dataf => N_31991,
datae => N_31998,
datad => N_31997,
datac => N_33264_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_30_RNIJN2QD_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_2\,
datae => N_32496,
datad => N_28580_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_24_3\(32),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff40")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_1\(30),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_334\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffccdc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_10\,
dataf => N_32903,
datae => N_32912,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datac => N_32278_2,
datab => N_32906,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_10_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff4000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_8\,
dataf => N_32914,
datae => N_32901,
datad => N_32925_2,
datac => N_31838_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_15_2_RNIBTVUH_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff80")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_11\,
dataf => N_32120,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_0\,
datad => N_32139,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datab => N_32135_2,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_1_RNI0JNF6_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff8000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_1\,
datae => N_33197,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(81),
datac => N_32221_1,
datab => N_32712_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffff2f02200")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_354\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2494\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2703\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2657\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffccdc0050")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_9\,
dataf => N_32983,
datae => N_31725_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_11_1\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_9_0\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0400")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2273\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1786\,
datad => N_27776_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(81),
datab => N_31715_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff20")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_4\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2609\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2582_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff20")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_11\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2274\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2697\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_1_22_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffff6f06600")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1071\,
dataf => N_33355,
datae => N_33001_1,
datad => N_33069,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2622_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_6_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffff0f1f1")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_318\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_6_3\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2652\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_6_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\(78));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_42: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0770088000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_42\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_25\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(39),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(38),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_40: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0078780000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_40\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_21\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_39: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0770088000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_39\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_19\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(49),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_38: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"14283c0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_38\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_17\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(43),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_46: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00003c0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_46\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_10\,
datae => N_79986,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_12\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_46_SUB: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fefbfdf7efbfdf7f")
port map (
combout => N_79986,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(19),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(11));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_COUNTSUCCESSIVEZERO36: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datad => N_79982,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_10\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_9\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_111_RNO_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"35ffffffffffffff")
port map (
combout => N_79935,
dataf => \GRLFPC2_0.FPO.FRAC\(49),
datae => \GRLFPC2_0.FPO.FRAC\(51),
datad => \GRLFPC2_0.FPO.FRAC\(47),
datac => N_26534,
datab => N_26574,
dataa => N_26573);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"569a569a569a66aa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10936\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10939\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"569a569a569a66aa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10935\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10939\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_26_RNIQV2S5_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333333337fffffff")
port map (
combout => N_79943,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2722\,
datae => N_31921_1,
datad => N_31766_2,
datac => N_31924_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_3_RNI8DAA6_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcccf000ffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2\,
dataf => N_79943,
datae => N_32619_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2776\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2490\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3_0\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_SUB_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfc0cfcfcfc0c0c0")
port map (
combout => N_79941,
dataf => N_28949,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742\,
datab => N_56);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_11_0_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff7f0000ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2466_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV\,
datae => N_79939,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_329\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN10_FEEDBACK\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_11_0_SUB_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"55ff55ff557f555f")
port map (
combout => N_79939,
dataf => N_79937,
datae => N_79923,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_329\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2757\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN10_FEEDBACK\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(73));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_110_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000707f0000f0ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV\,
datae => N_79937,
datad => N_79923,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN10_FEEDBACK\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(48));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN30_CONDITIONAL_0_RNIALVIO83: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"1090109010909090")
port map (
combout => N_79937,
dataf => \GRLFPC2_0.FPO.FRAC\(54),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN30_CONDITIONAL_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN10_FEEDBACK\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(48));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_111_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"2aaa2aaaeaaa2aaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT\(4),
dataf => N_79935,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_27_S_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(56));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_17_RNI6JB52: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00a200f700aa00ff")
port map (
combout => N_79923,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10920\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10918\,
datad => N_79931,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(50),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(49));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_21_RNI9AM21: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"a2a00200a0a20002")
port map (
combout => N_79931,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10924\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(50),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(49));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_17: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"faeefa4450ee5044")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10920\,
dataf => N_26592,
datae => N_26591,
datad => N_26534,
datac => N_26590,
datab => N_26589,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CHECKOVANDDENORM_UN13_NOTPOSSIBLEOV_5: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ca00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_5\,
dataf => \GRLFPC2_0.FPO.FRAC\(53),
datae => \GRLFPC2_0.FPO.FRAC\(52),
datad => \GRLFPC2_0.FPO.FRAC\(50),
datac => N_26534,
datab => N_26586,
dataa => N_26585);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_U: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000d0f00000505")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_2_2\,
datae => N_59229,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(42));
GRLFPC2_0_COMB_ANNULRES_1_IV: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff1110")
port map (
combout => \GRLFPC2_0.COMB.ANNULRES_1\,
dataf => \GRLFPC2_0.COMB.ANNULRES_1_IV_0\,
datae => \GRLFPC2_0.N_1676\,
datad => \GRLFPC2_0.ANNULRES_0_SQMUXA_10_0\,
datac => \GRLFPC2_0.N_1675_1\,
datab => \GRLFPC2_0.R.X.FPOP\,
dataa => \GRLFPC2_0.R.I.EXEC\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000009900f9f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_2\,
dataf => N_32739,
datae => N_32712_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_6_1\(25),
datac => N_31816_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O2_1_0_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fffcff000ffcc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O2_1\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c033000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_8\,
dataf => N_31725_1,
datae => N_32438_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O16_1_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f00000000000f00f")
port map (
combout => N_31983,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000fff000c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_9\,
dataf => N_33032,
datae => N_31775_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff4000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_9\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_0\,
datae => N_32852,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_19_1\(53),
datac => N_32786_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A12_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f020f0b0f000f000")
port map (
combout => N_33310,
dataf => N_31865_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(81),
datad => N_33333,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A12_0\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_49_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00aafcfc00aa0c0c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10093\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9797\,
datae => \GRLFPC2_0.FPI.LDOP_6\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(165),
dataa => N_700);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_9_0_RNIGCSSB_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"1505000011000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_10\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datae => N_32159,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccf0f0aaaaff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(55),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccaaaaf0f0ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(52),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccff00f0f0aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(48),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaff00ccccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(18),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_14_142_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0500ccccfa00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_14\(142),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(374),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(144),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(376));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0ccccff00aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(29),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccf0f0ff00aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(19),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_44_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaccccf0f0ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(44),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"e444a000a888a000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datae => N_33064_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2536\,
datac => N_32662_I,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ccccf0f0aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(32),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_42_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ccccf0f0aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(42),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaff00ccccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_41_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00aaaaf0f0cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(41),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ccccaaaaf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(8),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16));
GRLFPC2_0_V_FSR_AEXC_2_SQMUXA_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33f3ffffffffffff")
port map (
combout => \GRLFPC2_0.V.FSR.CEXC_3_SQMUXA_1\,
dataf => \GRLFPC2_0.N_1302\,
datae => \GRLFPC2_0.N_1720\,
datad => \GRLFPC2_0.COMB.ISFPOP2_1\,
datac => \GRLFPC2_0.R.X.LD\,
datab => \GRLFPC2_0.R.I.V\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffddddf0f0ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00cacaaa00aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7248\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4534\,
datae => \GRLFPC2_0.FPI.LDOP_4\,
datad => \GRLFPC2_0.FPI.OP1\(63),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3639\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(13));
GRLFPC2_0_R_A_RDD_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0f0f0f1f0")
port map (
combout => \GRLFPC2_0.R.A.RDD_0_0_G1\,
dataf => N_63,
datae => N_80,
datad => \GRLFPC2_0.COMB.RDD_1.M14_0_A2_3\,
datac => \GRLFPC2_0.N_73\,
datab => N_69,
dataa => N_59);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_3_0_0_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_3_0\(25),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_7_3_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000300000")
port map (
combout => N_32279_3,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_22_0_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_22_0\(52),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_A30_3_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0cfc000000000000")
port map (
combout => N_31922,
dataf => N_31886_2,
datae => N_32438_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_114_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000c000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(114),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(117));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_115_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000c000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(115),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(118));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_OPREXCSHFT_UN14_EXMIPTRLSBS_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffff000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2726\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(247),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(249),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(248));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_3_1_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000f00")
port map (
combout => N_32198_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_3_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3300cf0000000000")
port map (
combout => N_31713,
dataf => N_32272_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(81),
datad => N_31765_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_A26_3_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330000000f000000")
port map (
combout => N_32050,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(81),
datae => N_32050_1,
datad => N_31723_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A28_26_2_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000030fc0000")
port map (
combout => N_32413_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_O28_13_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff00ffffff00ff")
port map (
combout => N_32400,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O2_2_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c000ff00c000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O2_2\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_22_0_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f00000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_22_0\(57),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00030f0000030000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_12_TZ\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_9_1_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000f000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_9_1\(50),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_12_1_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2659\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_16_0_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f0000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_11_1\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_5_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f00000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2538\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_2_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3f30000000000000")
port map (
combout => N_32983,
dataf => N_32340_1,
datae => N_32434_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_6_1_44_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2622_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_3_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000c00000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2551\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_0_0_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c0000c0c00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A12_0_0\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_13_0_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f000f000f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_13_0\(36),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_1_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2490\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_2_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2498\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_A3_0_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2536\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_6_1_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_6_1\(25),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_15_0_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000300030000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_15_0\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A3_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2636\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_6_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000f00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2526\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_1_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"003f000000000000")
port map (
combout => N_31810,
dataf => N_31725_1_0,
datae => N_32120_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83),
datab => N_32048_1_0);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_2_2_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000ff")
port map (
combout => N_31811_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_13_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2268\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2671\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_18_RNIDBPB9_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff03000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_2\,
dataf => N_32484,
datae => N_32498_4,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_1_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f00000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2_1\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_1_0_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000000030f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A24_1_0\(33),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_O28_15_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff00ff00ff00")
port map (
combout => N_32404,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O2_1_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffcf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1164\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_10_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000300")
port map (
combout => N_33206,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_12_2_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f000000")
port map (
combout => N_32278_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_12_1_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000ff0000")
port map (
combout => N_32207_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_22_1_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000ff0000")
port map (
combout => N_32217_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_26_1_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000ff")
port map (
combout => N_32221_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A3_0_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000f0000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A3_0\(26),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_4_2_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff0000ff00")
port map (
combout => N_32057_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_20_1_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_31_1\(48),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_6_2_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccccc0000c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_6_2\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A28_16_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000000000000000")
port map (
combout => N_33072,
dataf => N_33136_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_0_0_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0cc0000000c00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0_0\(34),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_3_0_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A9_3_0\(28),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A28_8_1_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00000000000000")
port map (
combout => N_33064_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_0_0_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000c00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_0_0\(17),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_11_1_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000000000000")
port map (
combout => N_33207_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A28_31_1_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000000")
port map (
combout => N_32418_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fccccffffcccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10935\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_1_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0f0000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10865\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_61_RNIJNI68: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2599\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_2_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2633\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_1_0_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0303000000330000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A24_1_0\(55),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_11_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c000f0000000000")
port map (
combout => N_32586,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_4_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2508\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_2_3_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000c0000000000")
port map (
combout => N_32839_3,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_19_1_0_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_19_1\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_6_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000ffff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2648\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_23_0_A2_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8994\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_247\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(81),
datad => N_32048_1_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_15_0_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_15_0\(58),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_1_0_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff000000")
port map (
combout => N_31925_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_10_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"003c000000000000")
port map (
combout => N_32698,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(81),
datae => N_32425_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_10_1_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000003c00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A24_10_1\(55),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_4_0_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000cc0000000c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4_0\(59),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_17_2_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000ff")
port map (
combout => N_32289_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_8_0_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000fc00000030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_8_0\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_O26_0_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_32023,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O20_12_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0f0f0ff0f0f0f0")
port map (
combout => N_32336,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_6_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f0000000")
port map (
combout => N_33333,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_33_2_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f00000000000")
port map (
combout => N_32500_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_19_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000c00000000")
port map (
combout => N_32139,
dataf => N_31766_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A27_0_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000f0")
port map (
combout => N_31921_3,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A28_8_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f300000000000000")
port map (
combout => N_33064,
dataf => N_33136_1,
datae => N_31766_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_14_1_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff0000000000")
port map (
combout => N_32995_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_15_2_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff0000000000")
port map (
combout => N_32135_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_3_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0030000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2776\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_18_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300000000000000")
port map (
combout => N_32999,
dataf => N_32841_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3300300033000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2288\,
dataf => N_32344_1,
datae => N_33001_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2490\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_X2_3_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ffff000000ffff")
port map (
combout => N_32322_I,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_20_0_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f0f000f00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_20_0\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_5_37_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2689\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_12_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000c000000")
port map (
combout => N_33268,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_12_3_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000f00000")
port map (
combout => N_32619_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_9_0_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_9_0\(62),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_3_4_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000f0")
port map (
combout => N_33314_4,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_22_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000c00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2674\,
dataf => N_27776_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O2_0_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffff3ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_729\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(81),
datae => N_31763_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_21_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => N_32922,
dataf => N_32203_1,
datae => N_32487_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_21_1_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2576_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O3_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff00ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_255\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_10_3_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f3f000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_10_3\(59),
dataf => N_32066_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_6_0_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000fff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_6_0\(52),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_A30_12_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000c0000000")
port map (
combout => N_31931,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_9_0_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f0f0f00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_9_0\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_A30_12_1_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff000000")
port map (
combout => N_31931_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000f000000000")
port map (
combout => N_31808,
dataf => N_31803,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_19_2_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000f00000")
port map (
combout => N_32785_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_18_2_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f0000000000000")
port map (
combout => N_32784_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_32_4_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000f000")
port map (
combout => N_32498_4,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_4_1_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ff00")
port map (
combout => N_32290_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_12_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000003000f00030")
port map (
combout => N_32587,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_18_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000ff0000")
port map (
combout => N_33372,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_2_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000300000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2658\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_4_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2693\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_7_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0003000000000000")
port map (
combout => N_33360,
dataf => N_32841_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_5_0_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000ff")
port map (
combout => N_32243,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_41_2_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000f000")
port map (
combout => N_32563_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_17_0_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A24_17_0\(55),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_24_2_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00000000000000")
port map (
combout => N_32925_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_22_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000030000")
port map (
combout => N_32710,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_320\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(81),
datad => N_31892,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A28_24_0_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A28_24_0\(60),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_11_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000f00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_4914_1_A2_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_24_3_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0003000000000000")
port map (
combout => N_32712_3,
dataf => N_31839_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_6_1_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_6_1\(58),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_4_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f000c00000000")
port map (
combout => N_32841,
dataf => N_32841_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_3_3_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000300000")
port map (
combout => N_32840_3,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_5_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c3000000000000")
port map (
combout => N_32906,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_8_2_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f000000f00000")
port map (
combout => N_33264_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_19_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0030000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2341\,
dataf => N_32340_1_0,
datae => N_32203_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_7_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2283\,
dataf => N_32340_1_0,
datae => N_32203_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_7_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2504\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_15_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000300000000000")
port map (
combout => N_33271,
dataf => N_32069_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_3_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000300000")
port map (
combout => N_33356,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(81),
datae => N_31718_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_22_1_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_22_1\(52),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_14_2_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000f0000000000")
port map (
combout => N_33141_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_A29_22_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0030000000000000")
port map (
combout => N_32641,
dataf => N_32066_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_9_0_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_4_0\(34),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_6_1_A2_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000c00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2784\,
dataf => N_32066_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(78));
GRLFPC2_0_COMB_RDD_1_M14_0_A2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00000000000000")
port map (
combout => \GRLFPC2_0.COMB.RDD_1.M14_0_A2_3\,
dataf => N_81,
datae => \GRLFPC2_0.N_94\,
datad => \GRLFPC2_0.N_40\,
datac => N_72,
datab => N_74);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_A26_7_0_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_A26_7_0\(11),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccf0f0ff00ff00")
port map (
combout => N_59163,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccff00f0f0f0f0")
port map (
combout => N_59164,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0ff00ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8_I\(57),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(12));
\GRLFPC2_0_R_A_RF1REN_RNO_0_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000c0000000000")
port map (
combout => \GRLFPC2_0.COMB.V.A.RF1REN_1_0_7636_I_1\,
dataf => N_81,
datae => N_80,
datad => N_71,
datac => N_70,
datab => N_74);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_0_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f0000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2655\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A12_0_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A12_0\(61),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79));
GRLFPC2_0_COMB_UN3_IUEXEC_I_A3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.N_178\,
dataf => \GRLFPC2_0.R.X.FPOP\,
datae => \GRLFPC2_0.R.I.EXEC\,
datad => \GRLFPC2_0.R.E.FPOP\,
datac => \GRLFPC2_0.R.M.FPOP\,
datab => \GRLFPC2_0.R.A.FPOP\);
GRLFPC2_0_COMB_FPDECODE_FPOP2_0_A2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000c0000000000")
port map (
combout => \GRLFPC2_0.N_620\,
dataf => \GRLFPC2_0.N_77\,
datae => N_69,
datad => N_71,
datac => N_70,
datab => N_73);
GRLFPC2_0_COMB_FPDECODE_FPOP3_0_A2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00000000000000")
port map (
combout => \GRLFPC2_0.N_884\,
dataf => \GRLFPC2_0.N_77\,
datae => N_69,
datad => N_71,
datac => N_70,
datab => N_73);
\GRLFPC2_0_R_A_SEQERR_RET_4_RNIH90O2_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cf00000000000000")
port map (
combout => \GRLFPC2_0.R.A.AFQ\,
dataf => \GRLFPC2_0.N_27\,
datae => \GRLFPC2_0.R.E.AFQ_RET_0_0_G1_5\,
datad => \GRLFPC2_0.R.E.AFQ_RET_0_0_G1_4\,
datac => \GRLFPC2_0.R.STATE_O\(0),
datab => \GRLFPC2_0.R.STATE_O\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_11_2_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000f000")
port map (
combout => N_32206_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_20_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000c")
port map (
combout => N_32708,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(81),
datae => N_31892,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_11_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00300000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_1\,
dataf => N_32200,
datae => N_28580_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(81),
datac => N_31813_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83));
\GRLFPC2_0_R_STATE_RNIVPL21_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0003000300000003")
port map (
combout => \GRLFPC2_0.N_939_I_0_A2_2\,
dataf => \GRLFPC2_0.R.STATE\(1),
datae => \GRLFPC2_0.R.STATE\(0),
datad => N_85,
datac => N_84,
datab => N_10);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A17_0_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A17_0\(13),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A25_1_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000ff0000")
port map (
combout => N_33134_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A28_36_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000c")
port map (
combout => N_32423,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(81),
datae => N_32390_I,
datad => N_31788,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A28_38_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000c0000000000")
port map (
combout => N_32425,
dataf => N_33138_1,
datae => N_32142_1,
datad => N_32425_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A28_41_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000c0c00")
port map (
combout => N_32428,
dataf => N_32739,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A3_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000f00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2654\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_16_1_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000f000000000")
port map (
combout => N_33143_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_1_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2663\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_5_0_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000000")
port map (
combout => N_33133_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80));
GRLFPC2_0_COMB_FPDECODE_RDD5_0_A2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f00000000")
port map (
combout => \GRLFPC2_0.N_925\,
dataf => \GRLFPC2_0.N_93\,
datae => N_62,
datad => N_63,
datac => N_59);
GRLFPC2_0_COMB_RDD_1_M14_0_O2_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff0f000000")
port map (
combout => \GRLFPC2_0.N_38\,
dataf => N_61,
datae => N_60,
datad => N_58,
datac => N_57);
GRLFPC2_0_MOV_2_SQMUXA_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000c000000")
port map (
combout => \GRLFPC2_0.MOV_2_SQMUXA_1\,
dataf => N_61,
datae => \GRLFPC2_0.N_3418\,
datad => N_58,
datac => N_57,
datab => N_60);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffc0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_1\,
dataf => N_31867,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_3_0\(18),
datad => N_32070_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
GRLFPC2_0_COMB_ISFPOP2_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0f0f0f0f0f0")
port map (
combout => \GRLFPC2_0.COMB.ISFPOP2_1\,
dataf => \GRLFPC2_0.R.X.FPOP\,
datae => \GRLFPC2_0.R.I.V\,
datad => \GRLFPC2_0.R.I.EXEC\,
datac => \GRLFPC2_0.R.I.INST\(19),
datab => N_345);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_14_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300000000000000")
port map (
combout => N_32702,
dataf => N_28580_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_34_2_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f00000000")
port map (
combout => N_32567_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_0_0_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff30000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_6_RNI2NR84_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff30000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_2\,
dataf => N_31716,
datae => N_31743,
datad => N_31718_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_10_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff0cfff3ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(10),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(47),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(46),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00fff3ff0cffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(11),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(45),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(46),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_12_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00fff3ff0cffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(12),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(44),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(45),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00fff3ff0cffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(18),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(38),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(39),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff0cfff3ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(33),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(24),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(23),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00fff3ff0cffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(34),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(22),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(23),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_35_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff0cfff3ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(35),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(22),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(21),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00fff3ff0cffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(36),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(20),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(21),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_37_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff0cfff3ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(37),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(20),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(19),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_38_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00fff3ff0cffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(38),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(18),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(19),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_39_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00fff3ff0cffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(39),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_45_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff0cfff3ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(45),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(12),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff0cfff3ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(8),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(49),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_9_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00fff3ff0cffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(9),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(47),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_A26_14_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000300000")
port map (
combout => N_32061,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_16_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000c0000000")
port map (
combout => N_32136,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(81),
datae => N_32136_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_0_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000c00")
port map (
combout => N_32901,
dataf => N_28580_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(81),
datad => N_31813_2,
datac => N_31769_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_1_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff000000fff00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10868\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_1_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10872\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_1_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10870\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPYBUS_2_9_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(9),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_27: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03ff30000c00c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_27\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(40),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(45),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_17_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00000000000000")
port map (
combout => N_32998,
dataf => N_32487_2,
datae => N_32705_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_3_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccfff000cc00f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(238),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(251));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_4_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00030000000000")
port map (
combout => N_33260,
dataf => N_32487_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(81),
datad => N_32566_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_10_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => N_31998,
dataf => N_31766_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_1_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f0000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2513\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_1_9_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1967_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_21_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => N_32141,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(81),
datae => N_31766_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_3_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cc0000000f000000")
port map (
combout => N_32691,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(81),
datae => N_32425_1,
datad => N_31941_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_1_0_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000f0000000000")
port map (
combout => N_33069,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_34_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00000000000000")
port map (
combout => N_32500,
dataf => N_28580_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(81),
datad => N_31766_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_39_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1932\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(81),
datae => N_31715_1,
datad => N_32048_1_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_19_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2274\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2498\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_12_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1957\,
dataf => N_27776_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(81),
datad => N_31941_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_35_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c0000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2063\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2498\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_8_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000f000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2666\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffc0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1922\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2499\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_8_2_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff0000000000")
port map (
combout => N_32344_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_23_2_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00000000000000")
port map (
combout => N_32345_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_5_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => N_33261,
dataf => N_31766_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(81),
datad => N_32069_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_0_1_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c00c0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A9_0_1\(28),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNICRQFHA1_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff00fcfcfcfc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0\(9),
dataf => N_26534,
datae => N_26590,
datad => N_26588,
datac => N_26589,
datab => N_26587);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f0000f0000000")
port map (
combout => N_52547,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(81),
datae => N_52547_TZ,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN18_XZXBUS_14_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc0c03f3f0000fff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN18_XZXBUS_14\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(14),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_3_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c00c000000000000")
port map (
combout => N_33259,
dataf => N_32142_1,
datae => N_32066_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(78));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_21: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03ff30000c00c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_21\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(50),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_9_0_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff00ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_9_0\(19),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_17: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03ff30000c00c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_17\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_19: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f3f00c03000c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_19\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(56),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_19_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000c0000000000")
port map (
combout => N_33275,
dataf => N_31766_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(81),
datad => N_32566_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_19_1_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ff00")
port map (
combout => N_33275_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_23: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f3f00c03000c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_23\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(41),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_4_0_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c3c3c3c00ffff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_25: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03ff30000c00c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_25\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(36),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(37),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_21_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000c3000000")
port map (
combout => N_32487,
dataf => N_32739,
datae => N_32487_2,
datad => N_32566_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffcc0c33f30000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(8),
dataf => N_59194,
datae => N_59193,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_O26_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff000000ff00ffff")
port map (
combout => N_32093,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_23_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000c0000000")
port map (
combout => N_32143,
dataf => N_32020,
datae => N_31774_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_8_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000c00000000000")
port map (
combout => N_31817,
dataf => N_32340_1_0,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_247\,
datad => N_31788,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_9_0_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00000000000000")
port map (
combout => N_32159,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A28_29_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c0ff000000000000")
port map (
combout => N_32416,
dataf => N_31839_1,
datae => N_32908_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A3_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2763\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_10_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2697\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_6_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000300000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2788\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_18_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => N_33274,
dataf => N_31940_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(81),
datad => N_33136_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_27_S: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN10_FEEDBACK\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(50),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(49));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACKMULXFF_UN6_FEEDBACK: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(50),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(49));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_UN10_SELECTEDMIPTR_I_0_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0fff3ffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_I_0_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(76));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_UN10_SELECTEDMIPTR_I_0_O2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff0fffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(76));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTABORTNULLEXC_0_O2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ffff00ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(76));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_2_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000f000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2634\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_12_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000c00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2707\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_20_1_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000c000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2582_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_5_30_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2422\,
dataf => N_32340_1_0,
datae => N_31715_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A3_2_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2762\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_3_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c0000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2767\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_0_15_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2652\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_0_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2485\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_3_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f0000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2499\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_I_10_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000cfffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_10\(31),
dataf => N_31926,
datae => N_31813_2,
datad => N_31769_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_9_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => N_33136,
dataf => N_33136_1,
datae => N_32673_I,
datad => N_33136_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A28_47_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000003000000000")
port map (
combout => N_32434,
dataf => N_32908_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A3_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0030000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2586\,
dataf => N_33138_1,
datae => N_32203_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_13_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000300000000")
port map (
combout => N_32994,
dataf => N_32705_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_A26_2_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f3000300000000")
port map (
combout => N_32049,
dataf => N_31989_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_12_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000033000000000")
port map (
combout => N_32700,
dataf => N_31839_1,
datae => N_33298,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_30_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300000030000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1982\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(81),
datae => N_31763_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_0_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f00000f000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2602\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2494\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A3_21_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0030000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2779\,
dataf => N_32340_1_0,
datae => N_32048_1_0,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_3_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2706\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83),
datad => N_32048_1_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_1_20_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000300000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1931\,
dataf => N_31725_1_0,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_247\,
datad => N_32048_1_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A3_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2546\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_5_1_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000ff0000")
port map (
combout => N_31816_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_24_3_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f000f300000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_24_3\(32),
dataf => N_32688_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_1_2_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff000000")
port map (
combout => N_33312_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_25_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000c0000000000")
port map (
combout => N_32347,
dataf => N_31919_1,
datae => N_31774_1,
datad => N_31989_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_11_RNI7C1V4_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0c00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_2\,
dataf => N_31725_1,
datae => N_32131,
datad => N_32142_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A21_0_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000c0000000ccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A21_0\(59),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_A26_5_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000003000000000")
port map (
combout => N_32052,
dataf => N_31766_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(81),
datad => N_31723_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3300000003030000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2765\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(71),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(74),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(63));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffff0003300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_7\,
dataf => N_32853,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_6_1\(53),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_1_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => N_32838,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(81),
datae => N_32705_1,
datad => N_31691_I,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_22_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1967\,
dataf => N_32141_1_0,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_11_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000c0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1956\,
dataf => N_32343_1,
datae => N_32050_1,
datad => N_32136_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_3_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffcffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_647\,
dataf => N_32340_1_0,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_13_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000003000003")
port map (
combout => N_33367,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_9_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000ff")
port map (
combout => N_33023,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A28_0_0_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A28_0_0\(60),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(78));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_SA_I_1_0_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff3c3c00003c3c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1_0_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(316),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(258));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_5_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2703\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_37_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f00000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2505\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_9_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2319\,
dataf => N_31808_1,
datae => N_32048_1_0,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_4_43_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2534\,
dataf => N_32141_1_0,
datae => N_32048_1_0,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A3_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c0000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2725\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(81),
datae => N_32050_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_6_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000c00000")
port map (
combout => N_32907,
dataf => N_33040,
datae => N_32530_I,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_A3_0_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cc0c0000cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_A3_0_1\,
dataf => N_32203_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(66));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A3_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2484\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_15_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f030000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2337\,
dataf => N_31919_1,
datae => N_31924_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_A3_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2525\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0c000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_15\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_8\,
datae => N_32405,
datad => N_32908_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_19_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00000000000000")
port map (
combout => N_32785,
dataf => N_32141_1_0,
datae => N_31941_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_0_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000c0000")
port map (
combout => N_33256,
dataf => N_27553_1,
datae => N_32048_1,
datad => N_31989_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_21_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00000000000000")
port map (
combout => N_33277,
dataf => N_32141_1_0,
datae => N_32142_1,
datad => N_33136_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_28_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000300000000")
port map (
combout => N_32350,
dataf => N_32550_1,
datae => N_31724_1,
datad => N_33040,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_A30_10_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0030000000000000")
port map (
combout => N_31929,
dataf => N_32739,
datae => N_31813_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A28_35_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0003000003000000")
port map (
combout => N_32422,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(81),
datae => N_33063_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80));
GRLFPC2_0_COMB_ANNULRES_1_IV_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000fc00")
port map (
combout => \GRLFPC2_0.ANNULRES_0_SQMUXA_10_0\,
dataf => \GRLFPC2_0.R.E.FPOP\,
datae => \GRLFPC2_0.R.M.FPOP\,
datad => \GRLFPC2_0.R.A.FPOP\,
datac => N_153,
datab => N_154);
GRLFPC2_0_R_A_FPOP_RNIE2QG: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000000")
port map (
combout => \GRLFPC2_0.COMB.V.E.FPOP_1\,
dataf => \GRLFPC2_0.R.A.FPOP\,
datae => N_153,
datad => N_154);
GRLFPC2_0_R_E_LD_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000000")
port map (
combout => \GRLFPC2_0.R.E.LD_0_0_G1\,
dataf => \GRLFPC2_0.R.A.LD\,
datae => N_153,
datad => N_154);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A28_39_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000300000000000")
port map (
combout => N_32426,
dataf => N_33138_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A28_40_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c300000000000000")
port map (
combout => N_32427,
dataf => N_32066_2,
datae => N_31989_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_2_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000c00000000")
port map (
combout => N_32903,
dataf => N_31725_1_0,
datae => N_31766_1,
datad => N_31762_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O28_1_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030cc300000ff00")
port map (
combout => N_32894,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_2_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300300000000000")
port map (
combout => N_33355,
dataf => N_32272_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(81),
datad => N_31941_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_4_2_RNI6GGU5_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0030000000c00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19\(45),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(81),
datae => N_31763_1,
datad => N_31813_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_21_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03000c0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2127\,
dataf => N_32203_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(81),
datad => N_31762_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_10_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300000030000000")
port map (
combout => N_32911,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(81),
datae => N_31941_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff03000c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_8\,
dataf => N_33357,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datad => N_32120_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_9_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30c0000000000000")
port map (
combout => N_31997,
dataf => N_31775_1,
datae => N_31940_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(81),
datac => N_33136_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_3_30_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000c00000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2420\,
dataf => N_32203_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(81),
datad => N_32069_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_9_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff0000ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2598\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_12_0_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff0000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_12_0\(57),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_A29_3_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000003000000000")
port map (
combout => N_32622,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(81),
datae => N_31892,
datad => N_31718_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_10_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000030000")
port map (
combout => N_32130,
dataf => N_32070_1,
datae => N_31774_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(81),
datac => N_33040,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_O21_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff000000ffff")
port map (
combout => N_32246,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_16_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000000000000000")
port map (
combout => N_33143,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(81),
datae => N_32050_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_17_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000000000000000")
port map (
combout => N_33144,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(81),
datae => N_32050_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_I_A30_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0c0000000c0000")
port map (
combout => N_31918,
dataf => N_32070_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(81),
datad => N_31899_I,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_8_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00000000000000")
port map (
combout => N_33167,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_7_2_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f000000")
port map (
combout => N_33145_4,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_4_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => N_33357,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(81),
datae => N_31941_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_18_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => N_32784,
dataf => N_31839_1,
datae => N_31941_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_11_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0333000000000000")
port map (
combout => N_32777,
dataf => N_32645_3,
datae => N_31941_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A28_19_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => N_33075,
dataf => N_32142_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_13_0_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_13_0\(59),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_4_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030300000000000")
port map (
combout => N_32124,
dataf => N_31725_1_0,
datae => N_33063_1,
datad => N_31718_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_A29_7_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cf00000000000000")
port map (
combout => N_32626,
dataf => N_28580_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(81),
datad => N_32047_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_6_1_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_6_1\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_9_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000003000000")
port map (
combout => N_32846,
dataf => N_32739,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_320\,
datad => N_33071_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_25_0_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_25_0\(27),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_A30_25_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000c00000000000")
port map (
combout => N_31944,
dataf => N_32070_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A28_11_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000000000000000")
port map (
combout => N_33067,
dataf => N_32032_I,
datae => N_27297_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_6_10_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2302\,
dataf => N_32050_1,
datae => N_31723_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_4_30_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2421\,
dataf => N_32141_1_0,
datae => N_31715_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_1_37_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2518\,
dataf => N_31813_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A28_24_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c0000000000000")
port map (
combout => N_33080,
dataf => N_32141_1,
datae => N_31765_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A3_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000f00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2657\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_23_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0030000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2609\,
dataf => N_31725_1_0,
datae => N_32136_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_8_35_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0030000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2407\,
dataf => N_32066_2,
datae => N_31989_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_9_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000c000000")
port map (
combout => N_32281,
dataf => N_32141_1_0,
datae => N_32064_1,
datad => N_33063_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_11_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000c000000000")
port map (
combout => N_32131,
dataf => N_32064_1,
datae => N_31769_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2367\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_339\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_10_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c03000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2370\,
dataf => N_32908_1,
datae => N_32048_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_2_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1811\,
dataf => N_31725_1_0,
datae => N_32064_1,
datad => N_31924_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_7_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2560\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_11_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0c0000000000000")
port map (
combout => N_32992,
dataf => N_32487_2,
datae => N_33076_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(81),
datac => N_32048_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_1_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000003000")
port map (
combout => N_32273,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(81),
datae => N_32712_1,
datad => N_33063_1,
datac => N_33176,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_20_1_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000ff")
port map (
combout => N_33001_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_6_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0030000000000000")
port map (
combout => N_31769,
dataf => N_32487_2,
datae => N_32142_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(81),
datac => N_31769_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_A30_2_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000030000003300")
port map (
combout => N_31921,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_247\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(81),
datad => N_31766_2,
datac => N_33298,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_18_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000300000000000")
port map (
combout => N_33145,
dataf => N_32064_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(81),
datad => N_31813_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_11_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000003000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2354\,
dataf => N_32438_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(81),
datad => N_32662_I,
datac => N_32048_1_0,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_36_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000c00000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2214\,
dataf => N_27297_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(81),
datad => N_32069_2,
datac => N_33136_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_1_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000030000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1940\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(81),
datae => N_32120_1,
datad => N_32048_1_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_4_10_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000030000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2300\,
dataf => N_32438_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(81),
datad => N_32120_1,
datac => N_31924_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000030000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2369\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(81),
datae => N_32120_1,
datad => N_32390_I,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_6_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f00000000030000")
port map (
combout => N_32126,
dataf => N_31996_1,
datae => N_32064_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(81),
datac => N_33232,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000300000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2359\,
dataf => N_27776_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(81),
datad => N_31813_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_10_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000003000000")
port map (
combout => N_32991,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(81),
datae => N_32705_1,
datad => N_31899_I,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_3_1_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000ff")
port map (
combout => N_32128_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_3_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000ff")
port map (
combout => N_32932,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_0_14_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000000000")
port map (
combout => N_52211,
dataf => N_27776_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(81),
datad => N_32120_1,
datac => N_31718_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_19_1_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ff00")
port map (
combout => N_32485_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_20_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => N_33276,
dataf => N_31725_1_0,
datae => N_32438_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_O28_0_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff00ff")
port map (
combout => N_33032,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_6_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0003000000000000")
port map (
combout => N_33202,
dataf => N_27553_1,
datae => N_32422_1,
datad => N_32530_I,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_A26_6_1_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000c00000c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_A26_6_1\(11),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_1_RNIN2GH: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f033ff330fcc00cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_12239\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(258));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIV2O7_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff00000f0f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10635\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_0_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333cccc0ff00ff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24));
GRLFPC2_0_COMB_ANNULFPU_1_U_0_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcfcfcff000000")
port map (
combout => \GRLFPC2_0.COMB.ANNULFPU_1_U_0_0\,
dataf => \GRLFPC2_0.R.E.FPOP\,
datae => \GRLFPC2_0.R.A.FPOP\,
datad => \GRLFPC2_0.N_1237\,
datac => N_222,
datab => N_223);
GRLFPC2_0_R_M_FPOP_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000000")
port map (
combout => \GRLFPC2_0.R.M.FPOP_0_0_G1\,
dataf => \GRLFPC2_0.R.E.FPOP\,
datae => N_222,
datad => N_223);
GRLFPC2_0_R_M_LD_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000000")
port map (
combout => \GRLFPC2_0.R.M.LD_0_0_G1\,
dataf => \GRLFPC2_0.R.E.LD\,
datae => N_222,
datad => N_223);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_14_2_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000ff0000")
port map (
combout => N_32134_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_5_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000300000000")
port map (
combout => N_31768,
dataf => N_27929_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_320\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A28_4_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000030000")
port map (
combout => N_33060,
dataf => N_31688,
datae => N_33040,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_11_RNIJGRB5_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff03000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1956\,
datae => N_32550_1,
datad => N_31769_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A28_49_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000c0000000")
port map (
combout => N_32436,
dataf => N_31688,
datae => N_31763_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A28_37_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000c00000")
port map (
combout => N_32424,
dataf => N_33136_1,
datae => N_28580_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_11_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c0000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2321\,
dataf => N_32340_1_0,
datae => N_31762_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_8_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f300000000000000")
port map (
combout => N_32909,
dataf => N_32141_1,
datae => N_32435_1,
datad => N_31813_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_6_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff000000f000")
port map (
combout => N_31887,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A28_45_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => N_32432,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(81),
datae => N_32047_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_11_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0030000000000000")
port map (
combout => N_32699,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(81),
datae => N_32425_1,
datad => N_32662_I,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN8_TEMP_U_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"88088000ff7ff777")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10560\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10553\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10554\,
datac => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_0_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff00ff03333cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN1_CCIN: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fff0fff3333ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7210\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_0_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000c000000000")
port map (
combout => N_33127,
dataf => N_31724_1,
datae => N_32066_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(78));
GRLFPC2_0_R_X_FPOP_RNINRLL: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0003000000000000")
port map (
combout => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
dataf => \GRLFPC2_0.R.X.FPOP\,
datae => N_9,
datad => N_361,
datac => N_360,
datab => N_10);
GRLFPC2_0_COMB_ANNULRES_1_IV_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffc00030000")
port map (
combout => \GRLFPC2_0.COMB.ANNULRES_1_IV_0\,
dataf => \GRLFPC2_0.COMB.UN1_R.I.V_1\,
datae => \GRLFPC2_0.R.X.SEQERR\,
datad => N_361,
datac => N_360,
datab => N_10);
GRLFPC2_0_R_X_FPOP_RNIAQIJ: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f00000000")
port map (
combout => \GRLFPC2_0.V.I.EXEC_0_SQMUXA\,
dataf => \GRLFPC2_0.R.X.FPOP\,
datae => N_361,
datad => N_360,
datac => N_10);
GRLFPC2_0_V_FSR_FTT_3_SQMUXA_I_O2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffff0ffffffff")
port map (
combout => \GRLFPC2_0.N_3422\,
dataf => \GRLFPC2_0.R.X.SEQERR\,
datae => N_361,
datad => N_360,
datac => N_10);
GRLFPC2_0_R_X_AFSR_RNI0Q3P: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0003000000000000")
port map (
combout => \GRLFPC2_0.N_1132\,
dataf => \GRLFPC2_0.R.X.LD\,
datae => \GRLFPC2_0.R.X.AFSR\,
datad => N_361,
datac => N_360,
datab => N_10);
GRLFPC2_0_WRADDR_0_SQMUXA: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000030000")
port map (
combout => \GRLFPC2_0.N_1243\,
dataf => \GRLFPC2_0.R.X.AFSR\,
datae => \GRLFPC2_0.R.X.LD\,
datad => N_361,
datac => N_360,
datab => N_10);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_14_172_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000003000000fc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_14\(172),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(374),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(376));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_T_3_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0f3ff00f0f0cf0")
port map (
combout => N_59283,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(374),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(375),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(377),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(376));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN12_SRTOSTICKY_3_RNINBRL: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c0c0c0c0c0c0c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN12_SRTOSTICKY_3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_14_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f0f0fff0f0f0f")
port map (
combout => N_59162,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_16_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0f0f0f000f0f0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SCTRL_NEW\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_0_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c3c3c3c00ffff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN3_INEXACT: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000030303")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4664\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_28: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0003000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_28\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_26\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_20\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f00000f3f00300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10937\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0fc00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10944\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(43),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7782_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_10_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff33f3cc0c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(10),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(10),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_44_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffcc0c33f30000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(44),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(43),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42));
GRLFPC2_0_V_FSR_FTT_1_SQMUXA_3_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3fff3f0000ff3f")
port map (
combout => \GRLFPC2_0.V.FSR.FTT_1_SQMUXA_1\,
dataf => \GRLFPC2_0.R.X.LD\,
datae => \GRLFPC2_0.R.X.AFSR\,
datad => \GRLFPC2_0.R.STATE\(0),
datac => \GRLFPC2_0.R.STATE\(1),
datab => \GRLFPC2_0.R.X.AFQ\);
GRLFPC2_0_COMB_V_STATE2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff000000")
port map (
combout => \GRLFPC2_0.N_1213\,
dataf => \GRLFPC2_0.R.STATE\(0),
datae => \GRLFPC2_0.R.STATE\(1),
datad => \GRLFPC2_0.R.X.AFQ\);
GRLFPC2_0_COMB_V_FSR_RD_1_SN_M2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fffffff00000000")
port map (
combout => \GRLFPC2_0.N_3027\,
dataf => N_7,
datae => N_397,
datad => N_396,
datac => N_395);
GRLFPC2_0_V_STATE_0_SQMUXA: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000000000000000")
port map (
combout => \GRLFPC2_0.N_1669\,
dataf => N_431,
datae => N_397,
datad => N_396,
datac => N_395);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_27_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c0000c0000000000")
port map (
combout => N_32549,
dataf => N_33076_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(81),
datad => N_31718_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_7_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00c00000000000")
port map (
combout => N_32908,
dataf => N_32203_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(81),
datad => N_32908_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_15_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300300000000000")
port map (
combout => N_32210,
dataf => N_32131_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(81),
datad => N_31767_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN50_ZERO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f33fffffffff0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6961\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN48_ZERO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f33ffffffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN54_ZERO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000f33")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIN0DJ_49_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0ccf0ccf0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_372__G1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN35_ZERO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fffffffffccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6583\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN33_ZERO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fffffffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN20_ZERO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fffffffffccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5771\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNI64VE_21_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ccf0ccf0ccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5452\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN18_ZERO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fffffffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN24_ZERO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000330f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN39_ZERO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000330f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_7_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1816\,
dataf => N_31819_1,
datae => N_32438_1,
datad => N_32048_1_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_1_46_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1937\,
dataf => N_31819_1,
datae => N_32136_2,
datad => N_31924_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_3_37_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2579\,
dataf => N_31819_1,
datae => N_32487_2,
datad => N_31924_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_21_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1922\,
dataf => N_31819_1,
datae => N_32136_2,
datad => N_32048_1_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_1_1_RNICKDE4_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2373\,
dataf => N_31819_1,
datae => N_31763_1,
datad => N_31723_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_13_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0030000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2291\,
dataf => N_31819_1,
datae => N_31766_1,
datad => N_31723_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_22_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2544\,
dataf => N_31819_1,
datae => N_31899_I,
datad => N_31924_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_6_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000c0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2114\,
dataf => N_31819_1,
datae => N_32131_1,
datad => N_32136_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_0_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9471\,
dataf => N_31819_1,
datae => N_32438_1,
datad => N_31813_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_14_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000c0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2292\,
dataf => N_31725_1_0,
datae => N_32203_1,
datad => N_31762_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_24_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1969\,
dataf => N_31725_1_0,
datae => N_31762_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datac => N_32048_1_0,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_6_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1815\,
dataf => N_31921_1_0,
datae => N_31762_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_1_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33003300f3f03300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_334\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(81),
datae => N_31762_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2546\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff000c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_2\,
dataf => N_32986,
datae => N_32142_1,
datad => N_32064_1,
datac => N_31766_2,
datab => N_31769_1);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN14_CONDITIONAL_RNI3KDO2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000333")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5088\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1919\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_529\,
datac => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_2_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"030000000f000000")
port map (
combout => N_32768,
dataf => N_31688,
datae => N_33071_1,
datad => N_31765_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(11),
dataf => N_59192,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_12_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fccccccc0ccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_27_S_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(50),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccfffff0cc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(6),
dataf => N_59191,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A3_39_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2572\,
dataf => N_32120_1,
datae => N_32048_1_0,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_15_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcffffff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_15\(47),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_10\(47),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(81),
datad => N_32908_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_12_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3f00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2355\,
dataf => N_31921_1_0,
datae => N_31766_2,
datad => N_31924_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_21_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000c00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2590\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(81),
datae => N_31762_1,
datad => N_32673_I,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datab => N_32048_1_0);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_5_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc30cc0003cf33ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10883\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff30ba0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_3_0\(25),
datad => N_31899_I,
datac => N_31767_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_48_RNIJLN5B_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffff8f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2306\,
datad => N_31725_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2042\,
datab => N_27776_2,
dataa => N_31941_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00003000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_11\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9079\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_247\,
datad => N_31808_1,
datac => N_32048_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00030000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_7\,
dataf => N_33080,
datae => N_32438_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(81),
datac => N_31892,
datab => N_33232);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(13),
dataf => N_59215,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33000000b3008000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_9\,
dataf => N_28591_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4_0\(59),
datad => N_31763_1,
datac => N_32015_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_0_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0000000f000c000")
port map (
combout => N_32195,
dataf => N_31688,
datae => N_32620_1,
datad => N_31864_1,
datac => N_32047_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_14_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000030000000")
port map (
combout => N_32209,
dataf => N_31688,
datae => N_32022_I,
datad => N_31723_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_2_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1941\,
dataf => N_31996_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(81),
datad => N_31762_1,
datac => N_32050_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A2_4_0_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_4_0\(4),
dataf => N_32340_1_0,
datae => N_31996_1,
datad => N_31762_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\(78));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc0ff00ff033cc")
port map (
combout => N_58639,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f3cc3f00fc33cf0")
port map (
combout => N_58828,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(114),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc33cf00f3cc3f0")
port map (
combout => N_58361,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03fcf30c30cf3fc0")
port map (
combout => N_58384,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30cf3fc003fcf30c")
port map (
combout => N_58407,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f3cc3f00fc33cf0")
port map (
combout => N_58430,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc33cf00f3cc3f0")
port map (
combout => N_58453,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc30f3c3cf0c3f0")
port map (
combout => N_58476,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0fc33c3cc3f0f0")
port map (
combout => N_58499,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03fc30cff30c3fc0")
port map (
combout => N_58522,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30cf03fc3fc0f30c")
port map (
combout => N_58545,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0fc33c3cc3f0f0")
port map (
combout => N_58568,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03fcf30c30cf3fc0")
port map (
combout => N_58684,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03fc30cff30c3fc0")
port map (
combout => N_57901,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30cf03fc3fc0f30c")
port map (
combout => N_57924,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0fc33c3cc3f0f0")
port map (
combout => N_57947,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0fc33c3cc3f0f0")
port map (
combout => N_57970,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0fc33c3cc3f0f0")
port map (
combout => N_57993,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0fc33c3cc3f0f0")
port map (
combout => N_58016,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0fc33c3cc3f0f0")
port map (
combout => N_58039,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f3c0fc3c3f03cf0")
port map (
combout => N_58062,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc33cf00f3cc3f0")
port map (
combout => N_58085,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc33cf00f3cc3f0")
port map (
combout => N_58108,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fccf00f33f0cc")
port map (
combout => N_58707,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03fcf30c30cf3fc0")
port map (
combout => N_58131,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f33f0cc330fccf0")
port map (
combout => N_58154,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30cf3fc003fcf30c")
port map (
combout => N_58177,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc33cf00f3cc3f0")
port map (
combout => N_58200,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03fcf30c30cf3fc0")
port map (
combout => N_58223,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fccf00f33f0cc")
port map (
combout => N_57579,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30cf3fc003fcf30c")
port map (
combout => N_57602,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc30f3c3cf0c3f0")
port map (
combout => N_57625,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03fc30cff30c3fc0")
port map (
combout => N_57648,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30cf03fc3fc0f30c")
port map (
combout => N_57671,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fccf00f33f0cc")
port map (
combout => N_58730,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03fc30cff30c3fc0")
port map (
combout => N_57694,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30cf03fc3fc0f30c")
port map (
combout => N_57717,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03fc30cff30c3fc0")
port map (
combout => N_57740,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc0ff00ff033cc")
port map (
combout => N_57763,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff033cc33cc0ff0")
port map (
combout => N_57786,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c0f0f3c3cf0f03c")
port map (
combout => N_57809,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f3c3c0ff03c3cf0")
port map (
combout => N_57832,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc0ff00ff033cc")
port map (
combout => N_57855,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc0ff00ff033cc")
port map (
combout => N_57878,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc0ff00ff033cc")
port map (
combout => N_58593,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fccf00f33f0cc")
port map (
combout => N_58753,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc0ff00ff033cc")
port map (
combout => N_58616,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc0ff00ff033cc")
port map (
combout => N_58668,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c0f0f3c3cf0f03c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fccf00f33f0cc")
port map (
combout => N_58246,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fccf00f33f0cc")
port map (
combout => N_58269,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30cf3fc003fcf30c")
port map (
combout => N_58292,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc33cf00f3cc3f0")
port map (
combout => N_58315,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc33cf00f3cc3f0")
port map (
combout => N_58338,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_12_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => N_31875,
dataf => N_32627_1,
datae => N_32272_2,
datad => N_33298,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_40_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffccf00000ccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(40),
dataf => N_59206,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_9_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccc0cc00c0c00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_9\,
dataf => N_31819_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_39_0\(54),
datad => N_32487_2,
datac => N_31941_1,
datab => N_32220_1);
\GRLFPC2_0_COMB_V_FSR_FCC_1_1_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc30ff00ff00ff00")
port map (
combout => \GRLFPC2_0.N_3219\,
dataf => \GRLFPC2_0.R.X.LD\,
datae => \GRLFPC2_0.R.X.AFSR\,
datad => CPO_CCZ(0),
datac => N_373,
datab => \GRLFPC2_0.N_1105\);
\GRLFPC2_0_COMB_V_FSR_FCC_1_1_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc30ff00ff00ff00")
port map (
combout => \GRLFPC2_0.N_3220\,
dataf => \GRLFPC2_0.R.X.LD\,
datae => \GRLFPC2_0.R.X.AFSR\,
datad => CPO_CCZ(1),
datac => N_374,
datab => \GRLFPC2_0.N_1105\);
GRLFPC2_0_V_FSR_AEXC_1_SQMUXA_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f000000000000")
port map (
combout => \GRLFPC2_0.V.FSR.CEXC_2_SQMUXA_0\,
dataf => \GRLFPC2_0.R.X.LD\,
datae => \GRLFPC2_0.R.X.AFSR\,
datad => \GRLFPC2_0.N_1517\,
datac => \GRLFPC2_0.N_1105\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_39_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2581\,
dataf => N_32141_1_0,
datae => N_32120_1,
datad => N_31924_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_6_35_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000c0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2405\,
dataf => N_31921_1_0,
datae => N_32662_I,
datad => N_31924_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333333330000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_47__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2722\,
datae => N_33001_1,
datad => N_32136_2,
datac => N_31924_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_42_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000c0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2342\,
dataf => N_31921_1_0,
datae => N_32136_2,
datad => N_31924_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_43_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2263\,
dataf => N_31921_1_0,
datae => N_31899_I,
datad => N_31924_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN2_NOTDECODEDUNIMP_2_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000c00000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1902\,
dataf => N_32032_I,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_247\,
datad => N_32120_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2645\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_1_15_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1788\,
dataf => N_32141_1_0,
datae => N_32136_2,
datad => N_32048_1_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN1_MIFROMINST: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0c00000c000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3942\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_237\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(63));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff3000ffff3300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748\,
datae => \GRLFPC2_0.FPI.LDOP_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_237\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_74_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccccccccc0cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7274\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_237\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(62));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000f000f333f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_237\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_329\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_PCTRL_1_CO0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000fcff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_237\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_PCTRL_1_SUM_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff0300fcff")
port map (
combout => N_28945,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_237\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77));
GRLFPC2_0_COMB_ANNULFPU_1_U_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffc30")
port map (
combout => \GRLFPC2_0.COMB.ANNULFPU_1\,
dataf => \GRLFPC2_0.COMB.ANNULFPU_1_U_0_0\,
datae => \GRLFPC2_0.N_1675_1\,
datad => \GRLFPC2_0.R.X.FPOP\,
datac => \GRLFPC2_0.R.X.SEQERR\,
datab => \GRLFPC2_0.N_1105\);
GRLFPC2_0_WRADDR_1_SQMUXA: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffcfffcfffcf")
port map (
combout => \GRLFPC2_0.WRADDR_1_SQMUXA\,
dataf => \GRLFPC2_0.COMB.UN1_R.I.V_1\,
datae => \GRLFPC2_0.R.I.V\,
datad => \GRLFPC2_0.R.X.AFSR\,
datac => \GRLFPC2_0.R.X.LD\,
datab => \GRLFPC2_0.N_1105\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_6_A2_0_A2_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9079\,
dataf => N_32032_I,
datae => N_32203_1,
datad => N_31762_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_15_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1786\,
dataf => N_32141_1_0,
datae => N_33043_I,
datad => N_31924_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_13_RNIA2E93_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffc0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1958\,
datae => N_32141_1,
datad => N_31763_1,
datac => N_31813_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_13_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cc00c00000000000")
port map (
combout => N_32133,
dataf => N_32708_2,
datae => N_31768_1,
datad => N_32688_1,
datac => N_33063_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_5_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"003c000000000000")
port map (
combout => N_31814,
dataf => N_32340_1_0,
datae => N_32120_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_38_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffccf00000ccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(38),
dataf => N_59172,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffecffa0ffccff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_2\,
dataf => N_31819_1,
datae => N_32343_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2370\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_4914_1_A2_0\,
datab => N_32785_2,
dataa => N_32048_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_0_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f300f00000000000")
port map (
combout => N_32688,
dataf => N_32032_I,
datae => N_31763_1,
datad => N_32688_1,
datac => N_32425_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffff1f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2587\,
datae => N_33271,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2576_1\,
datac => N_33268,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_247\,
dataa => N_31723_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_19_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000300")
port map (
combout => N_32485,
dataf => N_31999_1,
datae => N_31921_1_0,
datad => N_32688_1,
datac => N_33232,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00c00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_2_1\,
dataf => N_31864,
datae => N_32627_1,
datad => N_33298,
datac => N_31769_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff30303000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_15\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_9\,
datae => N_32586,
datad => N_32587,
datac => N_32908_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffff4fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_14\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_8\,
datae => N_32894,
datad => N_32911,
datac => N_32907,
datab => N_31718_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_7_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f03000000000")
port map (
combout => N_32279,
dataf => N_32124_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(81),
datad => N_31691_I,
datac => N_32136_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0c0f00000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1808\,
dataf => N_32141_1_0,
datae => N_31763_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2599\,
datac => N_32120_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A18_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccc0000000000000")
port map (
combout => N_31709,
dataf => N_28591_1,
datae => N_31763_1,
datad => N_32015_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_9_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f5ff0000c4ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_9\(11),
dataf => N_32020,
datae => N_32048,
datad => N_31819_2,
datac => N_31788,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_9_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"eeaaeca0aaaaa0a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_3\,
dataf => N_32032_I,
datae => N_31999_1,
datad => N_31775_1,
datac => N_31762_1,
datab => N_32705_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A28_0_0\(60));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff50100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_5\,
dataf => N_32909,
datae => N_31999_1,
datad => N_32705_1,
datac => N_31813_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccc0ccc0ccc00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_647\,
datae => N_32136_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_329\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2757\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(73));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_3_1_RNIJICJ2_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff000000ffc8c8c8")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_14\,
dataf => N_32020,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_15_TZ\,
datad => N_32128_1,
datac => N_31775_1,
datab => N_32221_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccfffff0cc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(26),
dataf => N_59185,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff3cc3c33cff00")
port map (
combout => N_58070,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"030cfcf3cf3f30c0")
port map (
combout => N_58093,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_15_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2796\,
dataf => N_32203_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(81),
datad => N_31762_1,
datac => N_32050_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_8_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000030000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2318\,
dataf => N_32340_1_0,
datae => N_31763_1,
datad => N_31762_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_39_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ffffccf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(39),
dataf => N_59199,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_18_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000c0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2273\,
dataf => N_33138_1,
datae => N_31924_1,
datad => N_31989_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN2_NOTDECODEDUNIMP_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1903\,
dataf => N_32203_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2525\,
datac => N_32050_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2645\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_3_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1812\,
dataf => N_32487_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(81),
datad => N_32050_1,
datac => N_32048_1_0,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffc0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2321\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2490\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datac => N_31762_1,
datab => N_32050_1);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_NOTPROP_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30f0cf0fffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.NOTPROP_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN25_NOTPROP\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SCLSBS_2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_10_RNIS38G4_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff30303000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_1\,
dataf => N_32130,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datad => N_31865_1,
datac => N_31808_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CHECKOVANDDENORM_UN13_NOTPOSSIBLEOV: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_5\,
datae => \GRLFPC2_0.FPO.FRAC\(47),
datad => \GRLFPC2_0.FPO.FRAC\(51),
datac => \GRLFPC2_0.FPO.FRAC\(49),
datab => \GRLFPC2_0.FPO.FRAC\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0003000f000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_13\,
dataf => N_32141_1,
datae => N_32563_2,
datad => N_31723_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_5_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030300000300000")
port map (
combout => N_32277,
dataf => N_32246,
datae => N_32141_1_0,
datad => N_32064_1,
datac => N_31723_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccfffff0cc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(36),
dataf => N_59206,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_58601,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03cf0c3ffc30f3c0")
port map (
combout => N_58692,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(114),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c3f03cff3c0fc30")
port map (
combout => N_58392,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03f3303ffc0ccfc0")
port map (
combout => N_58415,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"303f03f3cfc0fc0c")
port map (
combout => N_58438,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03cf0c3ffc30f3c0")
port map (
combout => N_58461,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c033fcff3fcc030")
port map (
combout => N_58484,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c3ff3c3cffc300")
port map (
combout => N_58507,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ffc33c3cc3ff00")
port map (
combout => N_58530,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0330fccff33f0cc0")
port map (
combout => N_58553,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3003cffc3ff3c00c")
port map (
combout => N_58576,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ffc33c3cc3ff00")
port map (
combout => N_57909,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03f3303ffc0ccfc0")
port map (
combout => N_58715,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0330fccff33f0cc0")
port map (
combout => N_57932,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3003cffc3ff3c00c")
port map (
combout => N_57955,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ffc33c3cc3ff00")
port map (
combout => N_57978,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ffc33c3cc3ff00")
port map (
combout => N_58001,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ffc33c3cc3ff00")
port map (
combout => N_58024,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ffc33c3cc3ff00")
port map (
combout => N_58047,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c3f03cff3c0fc30")
port map (
combout => N_58116,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c3f03cff3c0fc30")
port map (
combout => N_58139,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_58738,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03f3303ffc0ccfc0")
port map (
combout => N_58162,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f33330ff0ccccf0")
port map (
combout => N_58185,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"303f03f3cfc0fc0c")
port map (
combout => N_58208,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c3f03cff3c0fc30")
port map (
combout => N_58231,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03f3303ffc0ccfc0")
port map (
combout => N_57587,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_57610,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30033ff3cffcc00c")
port map (
combout => N_57633,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c3ff3c3cffc300")
port map (
combout => N_57656,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0330fccff33f0cc0")
port map (
combout => N_57679,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3003cffc3ff3c00c")
port map (
combout => N_57702,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_58761,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0330fccff33f0cc0")
port map (
combout => N_57725,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3003cffc3ff3c00c")
port map (
combout => N_57748,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0330fccff33f0cc0")
port map (
combout => N_57771,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_57794,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f33330ff0ccccf0")
port map (
combout => N_57817,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3003cffc3ff3c00c")
port map (
combout => N_57840,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0330fccff33f0cc0")
port map (
combout => N_57863,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_57886,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_58624,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_58254,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_58647,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_58672,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_58277,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_58300,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"303f03f3cfc0fc0c")
port map (
combout => N_58323,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c3f03cff3c0fc30")
port map (
combout => N_58346,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c3f03cff3c0fc30")
port map (
combout => N_58369,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffff8f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_13\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8695\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_4\,
datad => N_33138_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2369\,
datab => N_32487_2,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2485\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_45_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ffffccf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(45),
dataf => N_59186,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_2_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3f0f0f033000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_346\,
dataf => N_31925_1,
datae => N_32050_1,
datad => N_31723_1,
datac => N_31813_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_9_12_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2311\,
dataf => N_32340_1_0,
datae => N_32487_2,
datad => N_32131_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_10_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1819\,
dataf => N_31725_1_0,
datae => N_32131_1,
datad => N_32136_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_A29_1_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3303000000000000")
port map (
combout => N_32620,
dataf => N_32620_1,
datae => N_32131_1,
datad => N_32120_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffff04ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_11\,
dataf => N_32545,
datae => N_32550_1,
datad => N_32549,
datac => N_32124_2,
datab => N_33076_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_7_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000c000000000")
port map (
combout => N_32773,
dataf => N_32340_1,
datae => N_31996_1,
datad => N_32632_1,
datac => N_32435_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_46_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(46),
dataf => N_59209,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_23_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccfffff0cc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(23),
dataf => N_59166,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_43_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(43),
dataf => N_59199,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccfffff0cc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(47),
dataf => N_59187,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_1_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"003c000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1810\,
dataf => N_32340_1_0,
datae => N_33064_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff30000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_568\,
datae => N_32340_1,
datad => N_32487_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2490\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(28),
dataf => N_59171,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_0_37_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffff444f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1042\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2579\,
datae => N_31921_1_0,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2655\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2499\,
datab => N_32784_2,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A25_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000300030000000")
port map (
combout => N_33126,
dataf => N_31775_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(81),
datad => N_32705_1,
datac => N_32047_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffccf00000ccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(51),
dataf => N_59187,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000c4c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_0\,
dataf => N_31865,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_320\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datac => N_32052_1,
datab => N_31769_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_37_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(37),
dataf => N_59180,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_49_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff4000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_7\,
dataf => N_32347,
datae => N_32357,
datad => N_31839_1,
datac => N_32705_1,
datab => N_32322_I,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff3000ffff2000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_4\,
dataf => N_32343_1,
datae => N_32998,
datad => N_31766_2,
datac => N_32220_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccfffff0cc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(33),
dataf => N_59180,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffff08ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_12\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_5\,
datae => N_28591_1,
datad => N_32848,
datac => N_31763_1,
datab => N_31762_1,
dataa => N_32908_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ffffccf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(25),
dataf => N_59174,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_3_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000003fffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_3\(11),
dataf => N_32061,
datae => N_32069_2,
datad => N_31819_2,
datac => N_32015_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_14_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000135f000033ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_14\(11),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_22_1\(52),
datae => N_32056,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_A26_7_0\(11),
datac => N_32390_I,
datab => N_32023,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_0_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ffffccf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(56),
dataf => N_59196,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff30c0ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_0\,
dataf => N_32141_1,
datae => N_32422,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83),
datac => N_32140_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_58615,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33333cc3c33ccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(114),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333c33c3cc3cccc")
port map (
combout => N_58337,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f3c3c0ff03c3cf0")
port map (
combout => N_58360,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c0f0f3c3cf0f03c")
port map (
combout => N_58383,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33333cc3c33ccccc")
port map (
combout => N_58406,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333c33c3cc3cccc")
port map (
combout => N_58429,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333c33c3cc3cccc")
port map (
combout => N_58452,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333c33c3cc3cccc")
port map (
combout => N_58475,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f3c3c0ff03c3cf0")
port map (
combout => N_58498,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c0f0f3c3cf0f03c")
port map (
combout => N_58521,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333c33c3cc3cccc")
port map (
combout => N_58544,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f3c3c0ff03c3cf0")
port map (
combout => N_58827,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f3c3c0ff03c3cf0")
port map (
combout => N_58567,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c0f0f3c3cf0f03c")
port map (
combout => N_57900,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333c33c3cc3cccc")
port map (
combout => N_57923,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333c33c3cc3cccc")
port map (
combout => N_57946,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333c33c3cc3cccc")
port map (
combout => N_57969,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333c33c3cc3cccc")
port map (
combout => N_57992,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333c33c3cc3cccc")
port map (
combout => N_58015,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333c33c3c3cc3ccc")
port map (
combout => N_58038,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33c33ccc333cc3cc")
port map (
combout => N_58061,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33c33ccc333cc3cc")
port map (
combout => N_58084,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc0ff00ff033cc")
port map (
combout => N_58683,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f3cf03c3c0f3cf0")
port map (
combout => N_58107,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff033cc33cc0ff0")
port map (
combout => N_58130,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c0f3cf00f3cf03c")
port map (
combout => N_58153,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33c33ccc333cc3cc")
port map (
combout => N_58176,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f3cf03c3c0f3cf0")
port map (
combout => N_58199,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc0ff00ff033cc")
port map (
combout => N_58222,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c0f0f3c3cf0f03c")
port map (
combout => N_57578,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333c33c3cc3cccc")
port map (
combout => N_57601,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f3c3c0ff03c3cf0")
port map (
combout => N_57624,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c0f0f3c3cf0f03c")
port map (
combout => N_57647,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc0ff00ff033cc")
port map (
combout => N_58706,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f3c3c0ff03c3cf0")
port map (
combout => N_57670,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c0f0f3c3cf0f03c")
port map (
combout => N_57693,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f3c3c0ff03c3cf0")
port map (
combout => N_57716,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_57739,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f33330ff0ccccf0")
port map (
combout => N_57762,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3003cffc3ff3c00c")
port map (
combout => N_57785,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0330fccff33f0cc0")
port map (
combout => N_57808,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_57831,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_57854,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_57877,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc0ff00ff033cc")
port map (
combout => N_58729,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_58592,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_58638,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3003cffc3ff3c00c")
port map (
combout => N_58667,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0330fccff33f0cc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc0ff00ff033cc")
port map (
combout => N_58752,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc0ff00ff033cc")
port map (
combout => N_58245,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c0f0f3c3cf0f03c")
port map (
combout => N_58268,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333c33c3cc3cccc")
port map (
combout => N_58291,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333c33c3cc3cccc")
port map (
combout => N_58314,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff80ffffff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_10\,
dataf => N_32032_I,
datae => N_33259,
datad => N_33271,
datac => N_32566_1,
datab => N_33136_2,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff9180ffff1100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_6\,
dataf => N_31886_2,
datae => N_32279,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_13_0\(59),
datac => N_32124_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff8f0ffff8800")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_13\,
dataf => N_33133_1,
datae => N_33126,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_5_2\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_6_0\(52),
datab => N_32908_1,
dataa => N_31768_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffc0ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_2\,
datae => N_31919_1,
datad => N_31989,
datac => N_32057_2,
datab => N_31989_1);
GRLFPC2_0_R_I_RDD_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000fc30ff00")
port map (
combout => \GRLFPC2_0.R.I.RDD_0_0_G1\,
dataf => \GRLFPC2_0.N_1470\,
datae => \GRLFPC2_0.R.X.FPOP\,
datad => \GRLFPC2_0.R.I.RDD\,
datac => \GRLFPC2_0.R.X.RDD\,
datab => \GRLFPC2_0.N_1105\);
GRLFPC2_0_V_FSR_FTT_3_SQMUXA_I_A3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0f0000ff000000")
port map (
combout => \GRLFPC2_0.V.FSR.FTT_3_SQMUXA_I_A3_0\,
dataf => \GRLFPC2_0.R.X.FPOP\,
datae => \GRLFPC2_0.R.I.V\,
datad => \GRLFPC2_0.R.I.EXEC\,
datac => \GRLFPC2_0.N_1105\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3f0f0f033000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_5\,
dataf => N_33264_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A24_1_0\(33),
datad => N_31766_1,
datac => N_33057_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A23_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3033000000000000")
port map (
combout => N_32980,
dataf => N_31725_1_0,
datae => N_31996_1,
datad => N_33232,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffff0f20022")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_7\,
dataf => N_32999,
datae => N_28591_1,
datad => N_32020,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_7_1\(6),
datab => N_32136_2,
dataa => N_31769_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_4_RNIEJT53_10_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00c00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_16__G2_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2300\,
datae => N_33133_1,
datad => N_31819_2,
datac => N_31723_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83));
\GRLFPC2_0_R_A_RF2REN_RNO_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0100030001000100")
port map (
combout => N_36381,
dataf => \GRLFPC2_0.N_178\,
datae => \GRLFPC2_0.N_1093\,
datad => N_81,
datac => N_80,
datab => N_36334,
dataa => \GRLFPC2_0.COMB.V.A.RF2REN_1_0_7690_I_A5_0_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_16\,
dataf => N_33256,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_5\,
datad => N_33277,
datac => N_32619_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_7_RNIJMS04_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffdc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_2\,
datae => N_33352,
datad => N_33360,
datac => N_33069,
datab => N_33357,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9074_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fefafcf0eeaacc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_2_0\,
dataf => N_31725_1,
datae => N_31921_3,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2788\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2526\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2508\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A3_0\(26));
\GRLFPC2_0_COMB_RS1_1_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcff30fffc003000")
port map (
combout => \GRLFPC2_0.COMB.RS1_1\(0),
dataf => \GRLFPC2_0.R.A.RS1\(0),
datae => N_64,
datad => N_9,
datac => \GRLFPC2_0.N_2989\,
datab => \GRLFPC2_0.N_889\);
\GRLFPC2_0_COMB_RS1_1_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcff30fffc003000")
port map (
combout => \GRLFPC2_0.COMB.RS1_1\(1),
dataf => \GRLFPC2_0.R.A.RS1\(1),
datae => N_65,
datad => N_9,
datac => \GRLFPC2_0.N_2990\,
datab => \GRLFPC2_0.N_889\);
\GRLFPC2_0_COMB_RS1_1_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcff30fffc003000")
port map (
combout => \GRLFPC2_0.COMB.RS1_1\(2),
dataf => \GRLFPC2_0.R.A.RS1\(2),
datae => N_66,
datad => N_9,
datac => \GRLFPC2_0.N_2991\,
datab => \GRLFPC2_0.N_889\);
\GRLFPC2_0_COMB_RS1_1_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcff30fffc003000")
port map (
combout => \GRLFPC2_0.COMB.RS1_1\(3),
dataf => \GRLFPC2_0.R.A.RS1\(3),
datae => N_67,
datad => N_9,
datac => \GRLFPC2_0.N_2992\,
datab => \GRLFPC2_0.N_889\);
\GRLFPC2_0_COMB_RS1_1_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcff30fffc003000")
port map (
combout => \GRLFPC2_0.COMB.RS1_1\(4),
dataf => \GRLFPC2_0.R.A.RS1\(4),
datae => N_68,
datad => N_9,
datac => \GRLFPC2_0.N_2993\,
datab => \GRLFPC2_0.N_889\);
\GRLFPC2_0_COMB_RS2_1_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ff00fff0000000")
port map (
combout => \GRLFPC2_0.COMB.RS2_1\(0),
dataf => \GRLFPC2_0.R.A.RS2\(0),
datae => N_50,
datad => N_9,
datac => \GRLFPC2_0.N_889\);
\GRLFPC2_0_COMB_RS2_1_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ff00fff0000000")
port map (
combout => \GRLFPC2_0.COMB.RS2_1\(1),
dataf => \GRLFPC2_0.R.A.RS2\(1),
datae => N_51,
datad => N_9,
datac => \GRLFPC2_0.N_889\);
\GRLFPC2_0_COMB_RS2_1_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ff00fff0000000")
port map (
combout => \GRLFPC2_0.COMB.RS2_1\(2),
dataf => \GRLFPC2_0.R.A.RS2\(2),
datae => N_52,
datad => N_9,
datac => \GRLFPC2_0.N_889\);
\GRLFPC2_0_COMB_RS2_1_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ff00fff0000000")
port map (
combout => \GRLFPC2_0.COMB.RS2_1\(3),
dataf => \GRLFPC2_0.R.A.RS2\(3),
datae => N_53,
datad => N_9,
datac => \GRLFPC2_0.N_889\);
\GRLFPC2_0_COMB_RS2_1_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ff00fff0000000")
port map (
combout => \GRLFPC2_0.COMB.RS2_1\(4),
dataf => \GRLFPC2_0.R.A.RS2\(4),
datae => N_54,
datad => N_9,
datac => \GRLFPC2_0.N_889\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_RNIMRL43_42_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff20")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_43__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_726\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_43__G2_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2342\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2508\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2484\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_RESULT_IV_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff05ff05ffcdff05")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\(12),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_I\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SFTLFT.AREGXORBREG_I_M\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN10_FEEDBACK\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(59));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_44_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_44__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_44__G2_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2534\,
datad => N_32619_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2490\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_24_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00f0f0ff00cccc")
port map (
combout => \GRLFPC2_0.N_3162\,
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.FSR.TEM\(1),
datac => N_687,
datab => N_623);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_21_RNIH7LP_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffc0ffffffea")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_255\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2674\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2590\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_339\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2490\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2582_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_O2_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffc0c0c0ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_354\,
dataf => N_33001_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2655\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2498\,
datac => N_32217_1,
datab => N_31723_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_1_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ffcc00f000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(13),
dataf => \GRLFPC2_0.FPI.OP2\(44),
datae => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_704,
datab => N_640);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_8_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc30cc0003cf33ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10886\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff3000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_12\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9074\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2373\,
datad => N_33133_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2634\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_46_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffccfcc33300300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(46),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(44),
datae => N_59209,
datad => N_59210,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_15_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(15),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(15),
datae => N_59215,
datad => N_59178,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_12_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bf370000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_12\(11),
dataf => N_31819_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_5\(11),
datad => N_33298,
datac => N_32057_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_MIFROMINST: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000cccccc0c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3924\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3942\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_255\,
datad => N_32136_2,
datac => N_33023,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.MIFROMINST_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff8")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_20\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_15\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_2\,
datac => N_33069,
datab => N_33032,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_6_1\(58));
\GRLFPC2_0_R_A_RF2REN_RNO_1_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000fff0")
port map (
combout => \GRLFPC2_0.COMB.V.A.RF2REN_1_0_7690_I_A5_0_0\,
dataf => N_82,
datae => N_83,
datad => \GRLFPC2_0.COMB.FPDECODE.ST\,
datac => \GRLFPC2_0.N_889\);
\GRLFPC2_0_COMB_V_E_STDATA_1_1_30_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00f0f0ff00cccc")
port map (
combout => \GRLFPC2_0.N_3168\,
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.FSR.RD\(0),
datac => N_693,
datab => N_629);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(13),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(13),
datae => N_59192,
datad => N_59173,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3ff333cc0cc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(28),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(28),
datae => N_59185,
datad => N_59220,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00f0f0ff00cccc")
port map (
combout => \GRLFPC2_0.N_3165\,
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.FSR.TEM\(4),
datac => N_690,
datab => N_626);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_12_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00c000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2290\,
dataf => N_33133_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2602\,
datad => N_32203_1,
datac => N_31762_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_24_RNINV1R1_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffc30cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_13\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1969\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2498\,
datad => N_32840_3,
datac => N_32120_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_1_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffecffa0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_1\(30),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2639\,
datae => N_32344_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2127\,
datac => N_32340_1_0,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2582_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2659\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_19_RNIEBLU7_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff84008800")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_4\,
dataf => N_32485,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_6_1\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
GRLFPC2_0_V_FSR_FTT_3_SQMUXA_I_O2_RNIDVU21: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffcc000f0f0c00")
port map (
combout => \GRLFPC2_0.N_1720\,
dataf => \GRLFPC2_0.N_1768\,
datae => \GRLFPC2_0.V.I.EXEC_0_SQMUXA\,
datad => \GRLFPC2_0.N_3422\,
datac => \GRLFPC2_0.R.I.V\,
datab => \GRLFPC2_0.R.I.EXEC\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff80")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_10\,
dataf => N_32287,
datae => N_32274,
datad => N_32280,
datac => N_32289_2,
datab => N_33071_1,
dataa => N_32140_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"eac0c0c0aa000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_11\,
dataf => N_31999_1,
datae => N_32932,
datad => N_32203_1,
datac => N_32632_1,
datab => N_33312_2,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_25_0\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_39_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffccfcc33300300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(39),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(37),
datae => N_59197,
datad => N_59199,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_1_22_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000030000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2640\,
dataf => N_27758_I,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2484\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffff8f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_18\,
dataf => N_32416,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_4\,
datad => N_33133_1,
datac => N_32421,
datab => N_32438_1,
dataa => N_32140_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_15_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffc0c0c0ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_596\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2494\,
datae => N_33143_1,
datad => N_31811_2,
datac => N_32048_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_0_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c0c00000ffc0ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_8__G2_0\,
dataf => N_31919_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2494\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2784\,
datac => N_32048_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_1_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ffccfff000cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(17),
dataf => \GRLFPC2_0.FPI.OP2\(37),
datae => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_703,
datab => N_639);
\GRLFPC2_0_COMB_V_E_STDATA_1_1_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00f0f0ff00cccc")
port map (
combout => \GRLFPC2_0.N_3163\,
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.FSR.TEM\(2),
datac => N_688,
datab => N_624);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffccfcc33300300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(25),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(23),
datae => N_59179,
datad => N_59174,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff8")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_14\,
dataf => N_33140,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_8\,
datad => N_33135,
datac => N_33127,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_7_0\(52),
dataa => N_33134_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffecff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2318\,
datae => N_32344_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2319\,
datac => N_31811_2,
datab => N_32840_3,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_885_I\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff80")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_3\,
datad => N_33355,
datac => N_32344_1,
datab => N_27297_1,
dataa => N_31941_1);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN1_CCIN_RNIJ2VG: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f03000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7035\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7210\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff80")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_11\,
dataf => N_32275,
datae => N_32272,
datad => N_32281,
datac => N_32290_1,
datab => N_32435_1,
dataa => N_31763_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_79_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ffcc00f000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(79),
dataf => \GRLFPC2_0.FPI.OP1\(36),
datae => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_664,
datab => N_600);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_82_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0ff00ccccff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(82),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => N_693,
datac => N_664,
datab => N_600);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_14_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3ff333cc0cc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(14),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(14),
datae => N_59183,
datad => N_59193,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00f0f0ff00cccc")
port map (
combout => \GRLFPC2_0.N_3144\,
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.FSR.AEXC\(1),
datac => N_669,
datab => N_605);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_68_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ffcc00f000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(68),
dataf => \GRLFPC2_0.FPI.OP1\(47),
datae => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_675,
datab => N_611);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_1_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ffccfff000cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(18),
dataf => \GRLFPC2_0.FPI.OP2\(36),
datae => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_702,
datab => N_638);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_RNI9IP62: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00c000c00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1281_I\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_2_1_CO1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_3_RNIL0F91: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00c000c00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_959_I\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_57\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_1_CO0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2_3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_3_RNIL0F91_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c0ff3fff3f00c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SBLSBS_2\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_57\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_1_CO0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2_3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_RNI19J12: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0fff0000f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_12247\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_2_1_CO1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_13_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_13\(11),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_4\(11),
datae => N_32052,
datad => N_32050);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_64_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ffccfff000cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(64),
dataf => \GRLFPC2_0.FPI.OP1\(48),
datae => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_682,
datab => N_618);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_40_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(40),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(40),
datae => N_59172,
datad => N_59208,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_63_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffc0ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1819\,
datae => N_32141_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1808\,
datac => N_31811_2,
datab => N_32048_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_83_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0ff00ccccff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(83),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => N_692,
datac => N_663,
datab => N_599);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffe000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_17\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_6\,
datad => N_32645_3,
datac => N_32142_1,
datab => N_31762_1,
dataa => N_32418_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_17\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_0\,
datae => N_32426,
datad => N_32428,
datac => N_32436,
datab => N_32423,
dataa => N_32434);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_63_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ffcc00f000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(63),
dataf => \GRLFPC2_0.FPI.OP1\(52),
datae => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_680,
datab => N_616);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff01010100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_0\,
datae => N_32141_1,
datad => N_33275_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_247\,
datab => N_32705_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3ff333cc0cc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(47),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(47),
datae => N_59186,
datad => N_59168,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
GRLFPC2_0_COMB_UN2_HOLDN_0_A3_7_RNIFSN01: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff80000000")
port map (
combout => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
dataf => \GRLFPC2_0.N_1255\,
datae => \GRLFPC2_0.COMB.UN2_HOLDN_0_A3_13\,
datad => \GRLFPC2_0.COMB.UN2_HOLDN_0_A3_11\,
datac => \GRLFPC2_0.COMB.UN2_HOLDN_0_A3_7\,
datab => \GRLFPC2_0.COMB.UN2_HOLDN_0_A3_10\,
dataa => \GRLFPC2_0.COMB.V.E.FPOP_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_60_Z_1_SUM_0_0_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c0ff3fff3f00c0")
port map (
combout => N_58671,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_12247\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2_3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_13\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2586\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2560\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_13_0\(36));
\GRLFPC2_0_R_E_STDATA_RNO_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"e400e4ffe400e400")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_28__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(60),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.R.I.PC\(28),
datab => \GRLFPC2_0.R.I.INST\(28),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_16_RNI1ELI5_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffff00ff40")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_6\,
dataf => N_32122,
datae => N_31921_1,
datad => N_32136,
datac => N_32134_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_23_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_23__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1071\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_23__G2_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1969\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2560\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2499\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_1_2_22_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffefacc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_1_2\(22),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2544\,
datae => N_32344_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2788\,
datac => N_32203_1,
datab => N_31763_1,
dataa => N_31931_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_6_RNI5466Q_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_17\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_7\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_1\,
datac => N_32126,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_10\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_14\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_1\,
datae => N_33261,
datad => N_33145_4,
datac => N_32142_1,
datab => N_33136_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_248_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffaa550030303030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(248),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10538\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10520\,
datad => \GRLFPC2_0.FPO.EXP\(9),
datac => \GRLFPC2_0.FPI.OP1\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_20_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3f00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_20\(11),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_9\(11),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_8\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_14\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1967_1\,
datab => N_32136_1);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN14_CONDITIONAL: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000033300000300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5088\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_6\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7144\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3848\,
datac => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233));
\GRLFPC2_0_R_E_STDATA_RNO_21_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"e400e4ffe400e400")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_21__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(53),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.R.I.PC\(21),
datab => \GRLFPC2_0.R.I.INST\(21),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A3_2_RNIGRHB2_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf0cc00f0f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_8\,
dataf => N_31725_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2513\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2505\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2762\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffff1fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_15\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_10\,
datae => N_31921_1,
datad => N_33275,
datac => N_33260,
datab => N_31788,
dataa => N_33232);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_30_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff80")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_30__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_1\(30),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_30__G2_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2422\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_334\,
datab => N_31924_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_24_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff8")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_24__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_1_2\(22),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_24__G2_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2640\,
datac => N_33355,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2513\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2657\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff8")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2291\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2292\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2663\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2538\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffeac0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_9\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_2_0\,
datad => N_32340_1,
datac => N_31725_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2706\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2659\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_16\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_10\,
datae => N_33148,
datad => N_33128,
datac => N_33144,
datab => N_33143);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffff888f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_10\,
dataf => N_32785,
datae => N_31839_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A24_1_0\(55),
datac => N_32066_2,
datab => N_32064_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A24_17_0\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"55045515ffaeffbf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(1),
dataf => N_59307,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8_I\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNITSA8_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
dataf => \GRLFPC2_0.FPI.LDOP_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datad => \GRLFPC2_0.R.MK.RST2\,
datac => N_7);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNISSA8_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000f000")
port map (
combout => N_76344,
dataf => \GRLFPC2_0.FPI.LDOP_1\,
datae => \GRLFPC2_0.R.MK.RST2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(5),
datac => N_7);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_68_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\,
dataf => \GRLFPC2_0.FPI.LDOP_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(12),
datad => \GRLFPC2_0.R.MK.RST2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(47),
datab => N_7);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_20\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_14\,
datae => N_52645,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_10\,
datac => N_32922);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O2_1_0_RNIU5EQ_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"030303030303030f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3729_I_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_318\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O2_2\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O2_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(66));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_30_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffcf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_30__G2_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2421\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2420\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2763\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2419\,
datab => N_31924_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3fcf0ff030c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(47),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(47),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(46),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff8")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_17\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_9\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_11\,
datad => N_32984,
datac => N_32992,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2655\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2498\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN2_MIXOIN_1_RNO_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f30c0cf30cf3f30c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5324\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5446\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(370));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_238_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffbf0000ff8c0000")
port map (
combout => N_36372,
dataf => \GRLFPC2_0.FPO.EXP\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_238__G2_0_7428_I_0\,
datad => \GRLFPC2_0.FPI.LDOP\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(251));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0f0f00ff3333")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(47),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffffff0f0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(51),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_242_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffbf0000ff8c0000")
port map (
combout => N_36368,
dataf => \GRLFPC2_0.FPO.EXP\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_242__G2_0_7304_I_0\,
datad => \GRLFPC2_0.FPI.LDOP\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(255));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_PCTRL_1_SUM_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ffff0003fcff00")
port map (
combout => N_28946,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3ccc3ccc33c33ccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10939\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10937\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ccf0ccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(11),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datae => N_59262,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_46_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0f0f00ff3333")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(46),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffffff0f0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(50),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_12_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000f0ccf0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(12),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datae => N_59258,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ccf0ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(31),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datae => N_59274,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_9\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_8\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2351\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2355\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffc00fcff0c000c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10129\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9833\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(13),
datad => \GRLFPC2_0.FPI.LDOP_6\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(129));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffc00fcff0c000c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10125\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9829\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(17),
datad => \GRLFPC2_0.FPI.LDOP_6\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(133));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffc00fcff0c000c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10124\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9828\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(18),
datad => \GRLFPC2_0.FPI.LDOP_6\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(134));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffff0ffff00f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10140\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9844\,
datae => \GRLFPC2_0.FPI.LDOP_6\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(118));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000fff0000000f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10087\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9791\,
datae => \GRLFPC2_0.FPI.LDOP_6\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(171));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000fff0000000f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10086\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9790\,
datae => \GRLFPC2_0.FPI.LDOP_6\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(172));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000fff0000000f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10085\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9789\,
datae => \GRLFPC2_0.FPI.LDOP_6\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(173));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_17\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_14\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_15\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_11\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_10\,
dataa => N_52474);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff33ffffff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(55),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(57),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"303000aafcfc00aa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10141\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.FPI.LDOP_6\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(117));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_240_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffbf0000ff8c0000")
port map (
combout => N_36370,
dataf => \GRLFPC2_0.FPO.EXP\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_240__G2_0_7366_I_0\,
datad => \GRLFPC2_0.FPI.LDOP\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(253));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_37_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0ccffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(37),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datae => N_59237,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000f0ccf0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(33),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datae => N_59237,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_23_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0ccffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(23),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datae => N_59272,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000f0ccf0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(27),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datae => N_59274,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff00ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(54),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0c00aafcfc00aa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10142\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.FPI.LDOP_6\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(116));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_243_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffbf0000ff8c0000")
port map (
combout => N_36367,
dataf => \GRLFPC2_0.FPO.EXP\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_243__G2_0_7273_I_0\,
datad => \GRLFPC2_0.FPI.LDOP\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(256));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_39_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0ccffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(39),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datae => N_59253,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_40_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ccf0ccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(40),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datae => N_59249,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_237_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffbf0000ff8c0000")
port map (
combout => N_36373,
dataf => \GRLFPC2_0.FPO.EXP\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_237__G2_0_7459_I_0\,
datad => \GRLFPC2_0.FPI.LDOP\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(250));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0f0fffff00ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(52),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0ccffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(26),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datae => N_59245,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_30_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000f0ccf0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(30),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datae => N_59242,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_A3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cccccccc000ccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2807\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5065\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_6\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3848\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNITL1C1_254_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffbf0000ff8c0000")
port map (
combout => N_36369,
dataf => \GRLFPC2_0.FPO.EXP\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_241__G2_0_7335_I_0\,
datad => \GRLFPC2_0.FPI.LDOP\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(254));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_45_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000f0ccf0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(45),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datae => N_59252,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff80")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_24\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_14\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_18\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_13\,
datac => N_32340_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2485\,
dataa => N_32066_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_239_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffbf0000ff8c0000")
port map (
combout => N_36371,
dataf => \GRLFPC2_0.FPO.EXP\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_239__G2_0_7397_I_0\,
datad => \GRLFPC2_0.FPI.LDOP\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(252));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_A3_RNIR5BR3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3729_I_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_A3_RNIIOM51: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3729_I_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422\,
datad => N_31762_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_A3_RNIKGEU2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M\(79),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3729_I_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_A3_RNILCEU2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M\(84),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3729_I_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742\);
GRLFPC2_0_COMB_V_FSR_FCC8: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000c0000000")
port map (
combout => \GRLFPC2_0.N_1515\,
dataf => \GRLFPC2_0.N_1721\,
datae => \GRLFPC2_0.N_1309\,
datad => \GRLFPC2_0.N_1720\,
datac => \GRLFPC2_0.COMB.ISFPOP2_1\,
datab => \GRLFPC2_0.R.I.V\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff00ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(56),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_63_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_4\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_6\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1816\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_568\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1815\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_244_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffbfff8c00000000")
port map (
combout => N_36366,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__G2_0_7242_I_0\,
datae => \GRLFPC2_0.FPO.EXP\(0),
datad => \GRLFPC2_0.FPI.LDOP\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(257));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ccf0ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(13),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datae => N_59265,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_21_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ccf0ccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(21),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datae => N_59234,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0ccffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(32),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datae => N_59240,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000f0ccf0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(36),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datae => N_59238,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_16_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ccf0ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(16),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datae => N_59258,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_20_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ccf0ccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(20),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datae => N_59260,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_22_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000f0ccf0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(22),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datae => N_59245,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ccf0ccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(18),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datae => N_59261,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ccf0ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(34),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datae => N_59242,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN2_MIXOIN_RNI64QJ1_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"030c0c3030c0c003")
port map (
combout => N_59287,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_947_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SALSBS_2\(0),
datad => N_59284,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SALSBS_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5446\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_12_RNIGI04I_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_11\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1967\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1957\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN14_CONDITIONAL_RNINBQC4: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000c000c0c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6_I\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5088\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2807\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_PCTRL_1_SUM_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3fffc000ffff0000")
port map (
combout => N_28949,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_PCTRL_1_CO3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_45_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0ccfffff0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(45),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(47),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datac => N_59252,
datab => N_59250);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_22_RNI7MFHI_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_9\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2674\,
datac => N_31743,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_1_TZ\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_39_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffccf00000ccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(39),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(41),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datac => N_59253,
datab => N_59254);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccfffff0cc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(31),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(31),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datac => N_59237,
datab => N_59236);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_21_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ffffccf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(21),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(21),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datac => N_59272,
datab => N_59273);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_40_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(40),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(42),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datac => N_59249,
datab => N_59238);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN2_NOTDECODEDUNIMP: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffaaff80ffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3926\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.STARTSHFT.UN2_NOTDECODEDUNIMP_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_445\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1903\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_334\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2485\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2645\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f00000033")
port map (
combout => N_59297,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ffffccf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(11),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(11),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datac => N_59265,
datab => N_59246);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcfffffffc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10205\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(55),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_20_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccfffff0cc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(20),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(20),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datac => N_59245,
datab => N_59261);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccfffff0cc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(34),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datac => N_59238,
datab => N_59243);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_71_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff000c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.UN36_PCTRL_NEW_I\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3924\,
datae => \GRLFPC2_0.N_1000\,
datad => \GRLFPC2_0.R.MK.RST\,
datac => \GRLFPC2_0.R.MK.RST2\,
datab => N_9);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_PCTRL_1_SUM_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff0f0f0f0f0f0f0")
port map (
combout => N_28950,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_PCTRL_1_SUM_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3cf0f0f0f0f0f0f0")
port map (
combout => N_28951,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23_1_SUM_0_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cc333cc33cc333cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1281_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_58\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7035\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7034\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_50_1_SUM_0_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cc333cc33cc333cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1281_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_58\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7035\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7051\);
GRLFPC2_0_COMB_V_I_EXEC_11_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000300")
port map (
combout => \GRLFPC2_0.COMB.V.I.EXEC_1_3\,
dataf => \GRLFPC2_0.N_1586\,
datae => \GRLFPC2_0.N_1515\,
datad => \GRLFPC2_0.N_1720\,
datac => \GRLFPC2_0.N_1470\,
datab => \GRLFPC2_0.COMB.ANNULRES_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30b8303074fc7474")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9789\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(115),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_TEMP: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00c0ffff00cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.TEMP\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748\,
datae => \GRLFPC2_0.FPI.LDOP_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(21));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_A3_RNIQDPF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cccc00c0cccc00cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748\,
datae => \GRLFPC2_0.FPI.LDOP_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIQM2H_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cccc00c0cccc00cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748\,
datae => \GRLFPC2_0.FPI.LDOP\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIG5SK4_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcfc0000fcfc00fc")
port map (
combout => N_76337,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6_I\,
datae => \GRLFPC2_0.FPI.LDOP_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_4_0_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c0c0c0cfc0c0cfc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_4_0\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742\,
datab => N_56);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_26_D: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fe32ef23dc10cd01")
port map (
combout => N_55054,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10920\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10924\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"5072d8fa5577ddff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(8),
dataf => N_59281,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_2_IV_RNO_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300330003000300")
port map (
combout => N_29788,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_I\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\,
datab => \GRLFPC2_0.FPI.LDOP_4\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNITT2I_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000fc00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10538\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\,
datad => \GRLFPC2_0.FPI.LDOP\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SS0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf0fc3000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4534\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897\,
datad => \GRLFPC2_0.FPI.LDOP\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2S2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3ffc30ff0f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4534\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897\,
datad => \GRLFPC2_0.FPI.LDOP\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_246_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00fff0f00000f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(246),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10536\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
datad => \GRLFPC2_0.FPI.LDOP_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_247_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30ff300030303030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(247),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10535\,
datad => \GRLFPC2_0.FPI.LDOP_4\,
datac => \GRLFPC2_0.FPI.OP1\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_249_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30ff300030303030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(249),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10533\,
datad => \GRLFPC2_0.FPI.LDOP_4\,
datac => \GRLFPC2_0.FPI.OP1\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_A29_5_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"9800320000000000")
port map (
combout => N_32624,
dataf => N_32131_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(81),
datad => N_32220_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_9_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff00")
port map (
combout => N_35958,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(21),
datae => \GRLFPC2_0.R.FSR.RD\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(1));
\GRLFPC2_0_COMB_DBGDATA_4_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3f3c0f3f3c0c0c0")
port map (
combout => CPO_DBG_DATAZ(7),
dataf => N_606,
datae => N_670,
datad => N_398,
datac => \GRLFPC2_0.R.FSR.AEXC\(2),
datab => N_397);
\GRLFPC2_0_COMB_DBGDATA_4_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3f3c0f3f3c0c0c0")
port map (
combout => CPO_DBG_DATAZ(8),
dataf => N_607,
datae => N_671,
datad => N_398,
datac => \GRLFPC2_0.R.FSR.AEXC\(3),
datab => N_397);
\GRLFPC2_0_COMB_DBGDATA_4_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3f3c0f3f3c0c0c0")
port map (
combout => CPO_DBG_DATAZ(11),
dataf => N_610,
datae => N_674,
datad => N_398,
datac => CPO_CCZ(1),
datab => N_397);
\GRLFPC2_0_COMB_DBGDATA_4_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3f3c0f3f3c0c0c0")
port map (
combout => CPO_DBG_DATAZ(5),
dataf => N_604,
datae => N_668,
datad => N_398,
datac => \GRLFPC2_0.R.FSR.AEXC\(0),
datab => N_397);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_5_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3202000000000000")
port map (
combout => N_32986,
dataf => N_31921_1_0,
datae => N_32136_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_4_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000200000000000")
port map (
combout => N_33131,
dataf => N_33138_1,
datae => N_32632_1,
datad => N_33232,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_4_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c0000080400000")
port map (
combout => N_32770,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(81),
datae => N_31941_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_8_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000e20000")
port map (
combout => N_33135,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_320\,
datae => N_31724_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_18_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0b01000000000000")
port map (
combout => N_32340,
dataf => N_32340_1,
datae => N_31838_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\(78));
\GRLFPC2_0_COMB_DBGDATA_4_10_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3f3c0f3f3c0c0c0")
port map (
combout => CPO_DBG_DATAZ(10),
dataf => N_609,
datae => N_673,
datad => N_398,
datac => CPO_CCZ(0),
datab => N_397);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A22_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000a800000")
port map (
combout => N_32836,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(81),
datae => N_32064_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\(78));
GRLFPC2_0_COMB_UN8_CCV_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff888f888f888")
port map (
combout => \GRLFPC2_0.COMB.UN8_CCV_2\,
dataf => N_207,
datae => \GRLFPC2_0.R.E.FPOP\,
datad => \GRLFPC2_0.R.X.FPOP\,
datac => N_345,
datab => \GRLFPC2_0.R.X.LD\,
dataa => \GRLFPC2_0.R.X.AFSR\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_1_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000020c000000000")
port map (
combout => N_33197,
dataf => N_33136_1,
datae => N_33040,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80));
GRLFPC2_0_COMB_V_A_SEQERR_1_0_O2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"008ac300008a008a")
port map (
combout => \GRLFPC2_0.N_10\,
dataf => \GRLFPC2_0.FPCI_O\(59),
datae => \GRLFPC2_0.FPCI_O\(58),
datad => \GRLFPC2_0.FPCI_O\(60),
datac => \GRLFPC2_0.R.STATE_O\(0),
datab => \GRLFPC2_0.R.STATE_O\(1),
dataa => \GRLFPC2_0.N_1837_O\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_2_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"a300000000000000")
port map (
combout => N_31865,
dataf => N_31865_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(81),
datad => N_31767_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\(78));
\GRLFPC2_0_COMB_DBGDATA_4_14_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3f3c0f3f3c0c0c0")
port map (
combout => CPO_DBG_DATAZ(14),
dataf => N_613,
datae => N_677,
datad => N_398,
datac => \GRLFPC2_0.R.FSR.FTT\(0),
datab => N_397);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_2_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"a0000000b0003000")
port map (
combout => N_32197,
dataf => N_32645_3,
datae => N_31766_1,
datad => N_32052_1,
datac => N_31941_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80));
GRLFPC2_0_R_FSR_NONSTD_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"b888b888fccc3000")
port map (
combout => \GRLFPC2_0.R.FSR.NONSTD_0_0_G1\,
dataf => \GRLFPC2_0.N_1132\,
datae => \GRLFPC2_0.R.FSR.NONSTD\,
datad => N_425,
datac => N_7,
datab => \GRLFPC2_0.N_3027\,
dataa => N_385);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_1_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000c000f0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9074\,
dataf => N_31921_1,
datae => N_32141_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9074_1\,
datac => N_31864_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_I_0_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"5f4c5f5fffccffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_0\(31),
dataf => N_32645_3,
datae => N_27553_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_320\,
datac => N_32422_1,
datab => N_31892,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A24_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c0c000000000000")
port map (
combout => N_32765,
dataf => N_31839_1,
datae => N_32015_1,
datad => N_32136_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_1_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c0c0000000c00000")
port map (
combout => N_33128,
dataf => N_32142_1,
datae => N_32124_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(81),
datac => N_32047_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M13_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0003000300030002")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M13\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_23_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"feeeeeeef0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_23__G2_0\,
dataf => N_33069,
datae => N_32217_1,
datad => N_31808_1,
datac => N_31723_1,
datab => N_31813_2,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_X2_1_RNI0VRPA_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffc0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_0\,
dataf => N_32497,
datae => N_28030_I,
datad => N_32052_1,
datac => N_31924_1,
datab => N_31989_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_RNITJED_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0033f0f30000f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_15_TZ\,
dataf => N_31996_1,
datae => N_31774_1,
datad => N_32064_1,
datac => N_31766_2,
datab => N_32434_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_3_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f000000330000")
port map (
combout => N_32984,
dataf => N_31725_1_0,
datae => N_32136_2,
datad => N_31788,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_2_RNIQBHB2_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff00ffc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_255\,
datae => N_32131_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2633\,
datac => N_32425_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A29_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"40cc404000000000")
port map (
combout => N_32194,
dataf => N_32141_1_0,
datae => N_32124_2,
datad => N_31763_1,
datac => N_32705_1,
datab => N_31941_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"44004400f4f04400")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_1\,
dataf => N_33136_1,
datae => N_32438_1,
datad => N_33071_1,
datac => N_33063_1,
datab => N_31765_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_4_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000c000000000")
port map (
combout => N_32985,
dataf => N_31921_1_0,
datae => N_32705_1,
datad => N_32566_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff4040ffff4000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_7\,
dataf => N_32141_1,
datae => N_32281,
datad => N_33138_1,
datac => N_32203_1,
datab => N_31775_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_39_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff400040004000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_39__G2_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2513\,
datae => N_27776_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2490\,
datac => N_32064_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(81),
dataa => N_32885_I);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_9_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bf838cb0bc808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10073\,
dataf => \GRLFPC2_0.FPO.FRAC\(47),
datae => \GRLFPC2_0.FPO.FRAC\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaa020000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_3\,
dataf => N_31921_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2498\,
datad => N_31763_1,
datac => N_31941_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_O2_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c0c00000d5c05500")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_445\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_255\,
datae => N_32340_1_0,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2525\,
datac => N_31763_1,
datab => N_31723_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_21_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3500000000000000")
port map (
combout => N_32343,
dataf => N_32343_1,
datae => N_32422_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\(78));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c0f3cf000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"6eeaf7bffb7f9dd5")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5301\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5339\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10888\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10890\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_18_2_RNI8PU55_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0303000057035500")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_2\,
dataf => N_31921_1,
datae => N_33207_1,
datad => N_32784_2,
datac => N_31899_I,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcccf000cccc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_3\,
dataf => N_31725_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2513\,
datad => N_32487_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2485\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2599\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0000000fc00cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_0\,
dataf => N_32739,
datae => N_32627_1,
datad => N_33076_1,
datac => N_32066_2,
datab => N_32069_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffc000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_4\,
dataf => N_33136_1,
datae => N_32210,
datad => N_32070_1,
datac => N_32435_1,
datab => N_33136_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f300c00033000000")
port map (
combout => N_52645,
dataf => N_32141_1,
datae => N_32032_I,
datad => N_32069_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_2_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000800")
port map (
combout => N_33129,
dataf => N_32142_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(81),
datad => N_32705_1,
datac => N_31768_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_38_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"b3a03300a0a00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2_0\,
dataf => N_32340_1,
datae => N_32345_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2498\,
datac => N_33043_I,
datab => N_32786_1,
dataa => N_32048_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_1_RNIAHIN3_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"dc50cc0050500000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_6_TZ\,
dataf => N_31921_1,
datae => N_32340_1,
datad => N_31766_1,
datac => N_28580_1,
datab => N_31838_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ae0c0c0caa000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_4\,
dataf => N_33001_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2494\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_320\,
datac => N_33043_I,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2652\,
dataa => N_31819_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_5_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c300000000000000")
port map (
combout => N_31993,
dataf => N_31921_1_0,
datae => N_32688_1,
datad => N_33136_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A28_2_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000c00")
port map (
combout => N_33058,
dataf => N_32438_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(81),
datad => N_31892,
datac => N_32566_1,
datab => N_31765_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f300000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_0\,
dataf => N_31688,
datae => N_31864_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_A29_2_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3300300000000000")
port map (
combout => N_32621,
dataf => N_32343_1,
datae => N_32066_2,
datad => N_31723_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0f0c0c000f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_0\,
dataf => N_31839_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_4_0\(34),
datad => N_33298,
datac => N_33040,
datab => N_32230);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M14S2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff00ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM12\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7782_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN11_WQSTSETS: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f7f7f707")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN11_WQSTSETS\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TEMP\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(14),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_0_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0003000f000000")
port map (
combout => N_32272,
dataf => N_28591_1,
datae => N_32141_1_0,
datad => N_32272_2,
datac => N_33232,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_2_1_RNI1RUE_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff000000ffc0c0c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_43__G2_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_255\,
datae => N_33001_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2498\,
datac => N_32136_2,
datab => N_32136_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_9_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000fc0000000000")
port map (
combout => N_31818,
dataf => N_32066_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(81),
datad => N_32159,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_10_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"eac0c0c0aa000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_0_1\,
dataf => N_32141_1,
datae => N_33138_1,
datad => N_31762_1,
datac => N_32705_1,
datab => N_31768_1,
dataa => N_31819_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_I_3_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cf45ff55cfcfffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_3\(31),
dataf => N_31839_1,
datae => N_32487_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_320\,
datac => N_32070_1,
datab => N_31788,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_49_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"88f8888800000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_4\,
dataf => N_32550_1,
datae => N_31724_1,
datad => N_32422_1,
datac => N_32705_1,
datab => N_31768_1,
dataa => N_31769_1);
\GRLFPC2_0_R_FSR_TEM_RNO_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"b888b888fccc3000")
port map (
combout => \GRLFPC2_0.R.FSR.TEM_1_0_2__G1\,
dataf => \GRLFPC2_0.N_1132\,
datae => \GRLFPC2_0.R.FSR.TEM\(2),
datad => N_428,
datac => N_7,
datab => \GRLFPC2_0.N_3027\,
dataa => N_388);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f4444444f0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_0\,
dataf => N_32032_I,
datae => N_27758_I,
datad => N_31996_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2654\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2_1\(5),
dataa => N_32022_I);
\GRLFPC2_0_R_FSR_TEM_RNO_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"b888b888fccc3000")
port map (
combout => \GRLFPC2_0.R.FSR.TEM_1_0_4__G1\,
dataf => \GRLFPC2_0.N_1132\,
datae => \GRLFPC2_0.R.FSR.TEM\(4),
datad => N_430,
datac => N_7,
datab => \GRLFPC2_0.N_3027\,
dataa => N_390);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_0_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"8000000010000000")
port map (
combout => N_31809,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(81),
datae => N_32712_1,
datad => N_32120_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\(78));
\GRLFPC2_0_R_FSR_RD_RNO_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"b888b888fccc3000")
port map (
combout => \GRLFPC2_0.R.FSR.RD_0_0_0__G1\,
dataf => \GRLFPC2_0.N_1132\,
datae => \GRLFPC2_0.R.FSR.RD\(0),
datad => N_433,
datac => N_7,
datab => \GRLFPC2_0.N_3027\,
dataa => N_393);
\GRLFPC2_0_R_FSR_RD_RNO_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"b888b888fccc3000")
port map (
combout => \GRLFPC2_0.R.FSR.RD_0_0_1__G1\,
dataf => \GRLFPC2_0.N_1132\,
datae => \GRLFPC2_0.R.FSR.RD\(1),
datad => N_434,
datac => N_7,
datab => \GRLFPC2_0.N_3027\,
dataa => N_394);
\GRLFPC2_0_R_FSR_TEM_RNO_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"b888b888fccc3000")
port map (
combout => \GRLFPC2_0.R.FSR.TEM_1_0_3__G1\,
dataf => \GRLFPC2_0.N_1132\,
datae => \GRLFPC2_0.R.FSR.TEM\(3),
datad => N_429,
datac => N_7,
datab => \GRLFPC2_0.N_3027\,
dataa => N_389);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_3_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000c000000000")
port map (
combout => N_31991,
dataf => N_32340_1_0,
datae => N_31940_1,
datad => N_32064_1,
datac => N_33063_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84));
\GRLFPC2_0_R_FSR_TEM_RNO_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"b888b888fccc3000")
port map (
combout => \GRLFPC2_0.R.FSR.TEM_1_0_1__G1\,
dataf => \GRLFPC2_0.N_1132\,
datae => \GRLFPC2_0.R.FSR.TEM\(1),
datad => N_427,
datac => N_7,
datab => \GRLFPC2_0.N_3027\,
dataa => N_387);
\GRLFPC2_0_R_FSR_TEM_RNO_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"b888b888fccc3000")
port map (
combout => \GRLFPC2_0.R.FSR.TEM_1_0_0__G1\,
dataf => \GRLFPC2_0.N_1132\,
datae => \GRLFPC2_0.R.FSR.TEM\(0),
datad => N_426,
datac => N_7,
datab => \GRLFPC2_0.N_3027\,
dataa => N_386);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0000000f000c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8639\,
dataf => N_32032_I,
datae => N_33133_1,
datad => N_32136_2,
datac => N_32136_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3373005000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_10\,
dataf => N_33167,
datae => N_32438_1,
datad => N_32050_1,
datac => N_31768_1,
datab => N_32047_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f030f0f0f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1954\,
dataf => N_32344_1,
datae => N_32995_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2654\,
datac => N_33023,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_1_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f004f0000004400")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2587\,
dataf => N_32925_2,
datae => N_27758_I,
datad => N_27297_1,
datac => N_32069_2,
datab => N_31723_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"5541414155000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_1\,
dataf => N_32708_2,
datae => N_32435_1,
datad => N_31989_1,
datac => N_33232,
datab => N_32645_2,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_6_RNIU5VP_10_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffecffa0ffccff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_16__G2_1\,
dataf => N_32340_1,
datae => N_32345_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2302\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2498\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2536\,
dataa => N_32662_I);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"dc505050cc000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_8\,
dataf => N_32645_3,
datae => N_33167,
datad => N_31724_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_6_1\(58),
datab => N_31808_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_34_RNI5BTJ5_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00220005")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_5_0\,
dataf => N_32500,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_247\,
datac => N_33232,
datab => N_33176,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_9_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff8f0ffff8800")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_3\,
dataf => N_32619_1,
datae => N_32500,
datad => N_33207_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2499\,
datab => N_31899_I,
dataa => N_31924_1);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c3c33cc00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(114),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_18_RNIVLJI3_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffc000c000c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_2\,
dataf => N_31921_1,
datae => N_33075,
datad => N_32066_2,
datac => N_33372,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffff8fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_9\,
dataf => N_32143,
datae => N_33133_1,
datad => N_33069,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8994\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_247\,
dataa => N_33063_1);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_6: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fda8dfdff7f72a7f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10872\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10887\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10885\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33));
\GRLFPC2_0_R_E_STDATA_RNO_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"44f044ff44f04400")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_1__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(33),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.R.FSR.CEXC\(1),
datab => \GRLFPC2_0.R.I.INST\(1),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cc000000fcf0f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_9\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_255\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2513\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2490\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2707\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_15_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_15__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2267\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_596\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1941\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1786\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1788\,
dataa => N_33145);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_243_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0ff000eeeeeeee")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_243__G2_0_7273_I_0\,
dataf => \GRLFPC2_0.FPI.LDOP\,
datae => \GRLFPC2_0.FPI.OP2\(53),
datad => \GRLFPC2_0.FPI.OP2\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_244_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0ff000eeeeeeee")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__G2_0_7242_I_0\,
dataf => \GRLFPC2_0.FPI.LDOP\,
datae => \GRLFPC2_0.FPI.OP2\(52),
datad => \GRLFPC2_0.FPI.OP2\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10));
\GRLFPC2_0_R_E_STDATA_RNO_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"44f044ff44f04400")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_0__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(32),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.R.FSR.CEXC\(0),
datab => \GRLFPC2_0.R.I.INST\(0),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_239_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0ff000eeeeeeee")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_239__G2_0_7397_I_0\,
dataf => \GRLFPC2_0.FPI.LDOP\,
datae => \GRLFPC2_0.FPI.OP2\(57),
datad => \GRLFPC2_0.FPI.OP2\(60),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffeca0fffffcf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_1\,
dataf => N_27758_I,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1982\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_9_1\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2526\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_9_0\(50),
dataa => N_32048_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_238_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0ff000eeeeeeee")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_238__G2_0_7428_I_0\,
dataf => \GRLFPC2_0.FPI.LDOP\,
datae => \GRLFPC2_0.FPI.OP2\(58),
datad => \GRLFPC2_0.FPI.OP2\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_35_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0cff000c0c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_35__G2_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2763\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2658\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2490\,
datac => N_32394_I,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_240_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0ff000eeeeeeee")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_240__G2_0_7366_I_0\,
dataf => \GRLFPC2_0.FPI.LDOP\,
datae => \GRLFPC2_0.FPI.OP2\(56),
datad => \GRLFPC2_0.FPI.OP2\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNI6I8I_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0ff000eeeeeeee")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_241__G2_0_7335_I_0\,
dataf => \GRLFPC2_0.FPI.LDOP\,
datae => \GRLFPC2_0.FPI.OP2\(55),
datad => \GRLFPC2_0.FPI.OP2\(58),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_237_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0ff000eeeeeeee")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_237__G2_0_7459_I_0\,
dataf => \GRLFPC2_0.FPI.LDOP\,
datae => \GRLFPC2_0.FPI.OP2\(59),
datad => \GRLFPC2_0.FPI.OP2\(62),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_242_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0ff000eeeeeeee")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_242__G2_0_7304_I_0\,
dataf => \GRLFPC2_0.FPI.LDOP\,
datae => \GRLFPC2_0.FPI.OP2\(54),
datad => \GRLFPC2_0.FPI.OP2\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f4f1f5fafefbff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(13),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(44),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(43),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f4f2f6f9fdfbff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(31),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(25),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(26),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(24),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_13: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ffc03fff00c03f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10916\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5088\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_44_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f8f2faf5fdf7ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(44),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(12),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f8f2faf5fdf7ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(17),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(39),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(40),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_14_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f9f4fdf2fbf6ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(14),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(43),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(41),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f9f4fdf2fbf6ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(56),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f1f4f5fafbfeff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(19),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(38),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(37),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_16_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f9f4fdf2fbf6ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(16),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(41),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(39),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(40),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_40_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f1f4f5fafbfeff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(40),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(15),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00000acc0acc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datae => N_59268,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000faccfacc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datae => N_59267,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f9f2fbf4fdf6ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(29),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(26),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(28),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_43_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f2f4f6f9fbfdff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(43),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(13),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(12),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(14),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_15_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f2f4f6f9fbfdff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(15),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(41),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(40),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f2f9fbf4f6fdff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(53),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_23_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f2f4f6f9fbfdff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(23),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(33),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_30_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f2f9fbf4f6fdff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(30),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(25),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(26),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_24_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f9f4fdf2fbf6ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(24),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(33),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_22_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f9f2fbf4fdf6ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(22),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(33),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(35),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccaaaaf0f0ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f8f2faf5fdf7ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(32),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(24),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(24),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_COMB_RF1REN_1_0_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f00dfd00f000f00")
port map (
combout => \GRLFPC2_0.N_3226\,
dataf => \GRLFPC2_0.N_889\,
datae => \GRLFPC2_0.COMB.LOCKGEN.LOCKI_I_I\,
datad => \GRLFPC2_0.R.A.RF1REN\(2),
datac => N_9,
datab => \GRLFPC2_0.COMB.RS2D_1\,
dataa => \GRLFPC2_0.COMB.RS2_1\(0));
\GRLFPC2_0_COMB_RF2REN_1_0_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfc0cfc0cfc00f00")
port map (
combout => \GRLFPC2_0.N_3033\,
dataf => \GRLFPC2_0.COMB.RS1_1\(0),
datae => \GRLFPC2_0.COMB.RS1D_1\,
datad => \GRLFPC2_0.R.A.RF2REN\(1),
datac => N_9,
datab => \GRLFPC2_0.COMB.V.A.RF2REN_1_1\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_BUSYMULXFF_UN2_TEMP_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"8888888000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.BUSYMULXFF.UN2_TEMP_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3926\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(70),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(68));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_9_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"50d872fa55dd77ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(9),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(9),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_245_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"afa0afa00000cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(245),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10538\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3639\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(245),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(232));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_250_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000fc30fc30")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(250),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10538\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10532\,
datad => \GRLFPC2_0.FPI.OP1\(62),
datac => \GRLFPC2_0.FPI.OP1\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_251_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcc3300f0f0f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(251),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10538\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10517\,
datad => \GRLFPC2_0.FPO.EXP\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_41\(251),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_252_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000fc30fc30")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(252),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10538\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10530\,
datad => \GRLFPC2_0.FPI.OP1\(60),
datac => \GRLFPC2_0.FPI.OP1\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_253_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000fc30fc30")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(253),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10538\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10529\,
datad => \GRLFPC2_0.FPI.OP1\(59),
datac => \GRLFPC2_0.FPI.OP1\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_254_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcc3300f0f0f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(254),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10538\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10514\,
datad => \GRLFPC2_0.FPO.EXP\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_41\(254),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_255_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcc3300f0f0f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(255),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10538\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10513\,
datad => \GRLFPC2_0.FPO.EXP\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_41\(255),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_256_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000f3c0f3c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(256),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10538\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10526\,
datad => \GRLFPC2_0.FPI.OP1\(53),
datac => \GRLFPC2_0.FPI.OP1\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_257_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000fc30fc30")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(257),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10538\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10525\,
datad => \GRLFPC2_0.FPI.OP1\(55),
datac => \GRLFPC2_0.FPI.OP1\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11));
\GRLFPC2_0_R_E_STDATA_RNO_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc30fffffc300000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_2__G1\,
dataf => \GRLFPC2_0.N_3140\,
datae => \GRLFPC2_0.R.A.AFQ\,
datad => \GRLFPC2_0.R.I.PC\(2),
datac => \GRLFPC2_0.R.I.INST\(2),
datab => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_R_E_STDATA_RNO_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc30fffffc300000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_3__G1\,
dataf => \GRLFPC2_0.N_3141\,
datae => \GRLFPC2_0.R.A.AFQ\,
datad => \GRLFPC2_0.R.I.PC\(3),
datac => \GRLFPC2_0.R.I.INST\(3),
datab => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_R_E_STDATA_RNO_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0fff0ccf000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_4__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(36),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_145\,
datab => \GRLFPC2_0.R.FSR.CEXC\(4));
\GRLFPC2_0_R_E_STDATA_RNO_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0fff0ccf000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_5__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(37),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_146\,
datab => \GRLFPC2_0.R.FSR.AEXC\(0));
\GRLFPC2_0_R_E_STDATA_RNO_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc30fffffc300000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_6__G1\,
dataf => \GRLFPC2_0.N_3144\,
datae => \GRLFPC2_0.R.A.AFQ\,
datad => \GRLFPC2_0.N_3426\,
datac => \GRLFPC2_0.R.I.INST\(6),
datab => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_R_E_STDATA_RNO_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc30fffffc300000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_7__G1\,
dataf => \GRLFPC2_0.N_3145\,
datae => \GRLFPC2_0.R.A.AFQ\,
datad => \GRLFPC2_0.N_3427\,
datac => \GRLFPC2_0.R.I.INST\(7),
datab => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_R_E_STDATA_RNO_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc30fffffc300000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_8__G1\,
dataf => \GRLFPC2_0.N_3146\,
datae => \GRLFPC2_0.R.A.AFQ\,
datad => \GRLFPC2_0.N_3428\,
datac => \GRLFPC2_0.R.I.INST\(8),
datab => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_R_E_STDATA_RNO_9_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc30fffffc300000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_9__G1\,
dataf => \GRLFPC2_0.N_3147\,
datae => \GRLFPC2_0.R.A.AFQ\,
datad => \GRLFPC2_0.N_3429\,
datac => \GRLFPC2_0.R.I.INST\(9),
datab => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_R_E_STDATA_RNO_10_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0fff0ccf000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_10__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(42),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_151\,
datab => CPO_CCZ(0));
\GRLFPC2_0_R_E_STDATA_RNO_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0fff0ccf000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_11__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(43),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_152\,
datab => CPO_CCZ(1));
\GRLFPC2_0_R_E_STDATA_RNO_12_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000f0fff000f000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_12__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(44),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_153\);
\GRLFPC2_0_R_E_STDATA_RNO_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc30fffffc300000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_13__G1\,
dataf => \GRLFPC2_0.N_3151\,
datae => \GRLFPC2_0.R.A.AFQ\,
datad => \GRLFPC2_0.N_140\,
datac => \GRLFPC2_0.R.I.INST\(13),
datab => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_R_E_STDATA_RNO_14_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc30fffffc300000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_14__G1\,
dataf => \GRLFPC2_0.N_3152\,
datae => \GRLFPC2_0.R.A.AFQ\,
datad => \GRLFPC2_0.N_141\,
datac => \GRLFPC2_0.R.I.INST\(14),
datab => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_R_E_STDATA_RNO_15_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000f0fff000f000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_15__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(47),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_156\);
\GRLFPC2_0_R_E_STDATA_RNO_16_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0fff0ccf000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_16__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(48),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_157\,
datab => \GRLFPC2_0.R.FSR.FTT\(2));
\GRLFPC2_0_R_E_STDATA_RNO_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0fff0fff0fff000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_17__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(49),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_3122\);
\GRLFPC2_0_R_E_STDATA_RNO_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc30fffffc300000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_18__G1\,
dataf => \GRLFPC2_0.N_3156\,
datae => \GRLFPC2_0.R.A.AFQ\,
datad => \GRLFPC2_0.R.I.PC\(18),
datac => \GRLFPC2_0.R.I.INST\(18),
datab => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_R_E_STDATA_RNO_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000f0fff000f000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_19__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(51),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_158\);
\GRLFPC2_0_R_E_STDATA_RNO_20_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000f0fff000f000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_20__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(52),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_3125\);
\GRLFPC2_0_R_E_STDATA_RNO_22_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc30fffffc300000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_22__G1\,
dataf => \GRLFPC2_0.N_3160\,
datae => \GRLFPC2_0.R.A.AFQ\,
datad => \GRLFPC2_0.R.I.PC\(22),
datac => \GRLFPC2_0.R.I.INST\(22),
datab => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_R_E_STDATA_RNO_23_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0fff0ccf000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_23__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(55),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_3128\,
datab => \GRLFPC2_0.R.FSR.TEM\(0));
\GRLFPC2_0_R_E_STDATA_RNO_24_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc30fffffc300000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_24__G1\,
dataf => \GRLFPC2_0.N_3162\,
datae => \GRLFPC2_0.R.A.AFQ\,
datad => \GRLFPC2_0.R.I.PC\(24),
datac => \GRLFPC2_0.R.I.INST\(24),
datab => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_R_E_STDATA_RNO_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc30fffffc300000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_25__G1\,
dataf => \GRLFPC2_0.N_3163\,
datae => \GRLFPC2_0.R.A.AFQ\,
datad => \GRLFPC2_0.R.I.PC\(25),
datac => \GRLFPC2_0.R.I.INST\(25),
datab => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_R_E_STDATA_RNO_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc30fffffc300000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_26__G1\,
dataf => \GRLFPC2_0.N_3164\,
datae => \GRLFPC2_0.R.A.AFQ\,
datad => \GRLFPC2_0.R.I.PC\(26),
datac => \GRLFPC2_0.R.I.INST\(26),
datab => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_R_E_STDATA_RNO_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc30fffffc300000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_27__G1\,
dataf => \GRLFPC2_0.N_3165\,
datae => \GRLFPC2_0.R.A.AFQ\,
datad => \GRLFPC2_0.R.I.PC\(27),
datac => \GRLFPC2_0.R.I.INST\(27),
datab => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_R_E_STDATA_RNO_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000f0fff000f000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_29__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(61),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_3134\);
\GRLFPC2_0_R_E_STDATA_RNO_30_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc30fffffc300000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_30__G1\,
dataf => \GRLFPC2_0.N_3168\,
datae => \GRLFPC2_0.R.A.AFQ\,
datad => \GRLFPC2_0.R.I.PC\(30),
datac => \GRLFPC2_0.R.I.INST\(30),
datab => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_R_E_STDATA_RNO_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0fff0ccf000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_31__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(63),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_3136\,
datab => \GRLFPC2_0.R.FSR.RD\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00fffcff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\,
datad => \GRLFPC2_0.FPI.LDOP_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPBREGLOADEN: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00fffcff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\,
datad => \GRLFPC2_0.FPI.LDOP_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25));
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_0_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfc0c0c0cfcfcfcf")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV_0\(0),
dataf => \GRLFPC2_0.N_1570\,
datae => \GRLFPC2_0.R.FSR.TEM\(0),
datad => \GRLFPC2_0.R.I.EXC\(0),
datac => \GRLFPC2_0.N_1517\,
datab => N_403);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_0_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfc0c0c0cfcfcfcf")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV_0\(1),
dataf => \GRLFPC2_0.N_1570\,
datae => \GRLFPC2_0.R.FSR.TEM\(1),
datad => \GRLFPC2_0.R.I.EXC\(1),
datac => \GRLFPC2_0.N_1517\,
datab => N_404);
GRLFPC2_0_V_STATE_0_SQMUXA_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00000000000000")
port map (
combout => \GRLFPC2_0.N_1517\,
dataf => N_395,
datae => N_396,
datad => N_397);
GRLFPC2_0_COMB_UN2_HOLDN_0_A3_8: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f000f000f")
port map (
combout => \GRLFPC2_0.COMB.UN2_HOLDN_0_A3_8\,
dataf => \GRLFPC2_0.FPCI_O\(47),
datae => \GRLFPC2_0.FPCI_O\(46),
datad => \GRLFPC2_0.FPCI_O\(51),
datac => \GRLFPC2_0.FPCI_O\(50));
GRLFPC2_0_COMB_UN2_HOLDN_0_A3_13: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000030000000000")
port map (
combout => \GRLFPC2_0.COMB.UN2_HOLDN_0_A3_13\,
dataf => \GRLFPC2_0.COMB.UN2_HOLDN_0_A3_8\,
datae => \GRLFPC2_0.FPCI_O\(49),
datad => \GRLFPC2_0.FPCI_O\(44),
datac => \GRLFPC2_0.FPCI_O\(48),
datab => \GRLFPC2_0.FPCI_O\(45));
GRLFPC2_0_COMB_UN2_HOLDN_0_A3_7: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => \GRLFPC2_0.COMB.UN2_HOLDN_0_A3_7\,
dataf => \GRLFPC2_0.FPCI_O\(62),
datae => \GRLFPC2_0.FPCI_O\(69));
GRLFPC2_0_COMB_UN2_HOLDN_0_A3_11: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000f00000")
port map (
combout => \GRLFPC2_0.COMB.UN2_HOLDN_0_A3_11\,
dataf => \GRLFPC2_0.FPCI_O\(59),
datae => \GRLFPC2_0.FPCI_O\(60),
datad => \GRLFPC2_0.FPCI_O\(58),
datac => \GRLFPC2_0.FPCI_O\(70));
GRLFPC2_0_COMB_UN2_HOLDN_0_A3_10: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000f000000000")
port map (
combout => \GRLFPC2_0.COMB.UN2_HOLDN_0_A3_10\,
dataf => \GRLFPC2_0.FPCI_O\(63),
datae => \GRLFPC2_0.FPCI_O\(61),
datad => \GRLFPC2_0.FPCI_O\(52),
datac => N_9);
GRLFPC2_0_COMB_UN8_CCV: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000003f3f3f")
port map (
combout => CPO_CCVZ,
dataf => \GRLFPC2_0.COMB.UN8_CCV_2\,
datae => \GRLFPC2_0.R.M.FPOP\,
datad => N_276,
datac => \GRLFPC2_0.R.I.INST\(19),
datab => \GRLFPC2_0.R.I.EXEC\);
\GRLFPC2_0_R_A_AFQ_RET_RNIPDCL_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f0000000")
port map (
combout => \GRLFPC2_0.R.E.AFQ_RET_0_0_G1_5\,
dataf => \GRLFPC2_0.FPCI_O\(62),
datae => \GRLFPC2_0.FPCI_O\(69),
datad => \GRLFPC2_0.FPCI_O\(59),
datac => \GRLFPC2_0.FPCI_O\(60));
\GRLFPC2_0_R_A_AFQ_RET_RNINCIR_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000f00000")
port map (
combout => \GRLFPC2_0.R.E.AFQ_RET_0_0_G1_4\,
dataf => \GRLFPC2_0.FPCI_O\(61),
datae => \GRLFPC2_0.FPCI_O\(63),
datad => \GRLFPC2_0.FPCI_O\(58),
datac => \GRLFPC2_0.FPCI_O\(70));
GRLFPC2_0_R_E_SEQERR_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00000000000000")
port map (
combout => \GRLFPC2_0.R.E.SEQERR_0_0_G1\,
dataf => \GRLFPC2_0.N_11\,
datae => \GRLFPC2_0.N_27\,
datad => \GRLFPC2_0.FPCI_O\(70),
datac => \GRLFPC2_0.FPCI_O\(61),
datab => \GRLFPC2_0.FPCI_O\(63));
\GRLFPC2_0_R_A_AFQ_RET_RNI069S_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000c00000")
port map (
combout => \GRLFPC2_0.R.E.AFSR_RET_0_0_G1_3\,
dataf => \GRLFPC2_0.FPCI_O\(62),
datae => \GRLFPC2_0.FPCI_O\(69),
datad => \GRLFPC2_0.FPCI_O\(59),
datac => \GRLFPC2_0.FPCI_O\(70),
datab => \GRLFPC2_0.FPCI_O\(58));
GRLFPC2_0_COMB_UN1_FPCI_3_1_0_O2_RNIMTJ72: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00000000000000")
port map (
combout => \GRLFPC2_0.R.A.AFSR\,
dataf => \GRLFPC2_0.N_27\,
datae => \GRLFPC2_0.R.E.AFSR_RET_0_0_G1_3\,
datad => \GRLFPC2_0.N_7\,
datac => \GRLFPC2_0.FPCI_O\(61),
datab => \GRLFPC2_0.FPCI_O\(63));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_2_RNI51QB6_0_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff30000003ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(374),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(0));
GRLFPC2_0_R_MK_BUSY2_RET_1_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f00000000000")
port map (
combout => \GRLFPC2_0.N_2111\,
dataf => \GRLFPC2_0.R.MK.BUSY_4\,
datae => \GRLFPC2_0.R.MK.RST_O_0\,
datad => \GRLFPC2_0.R.MK.HOLDN2_O_0\,
datac => N_7);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_0_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfc0c0c0cfcfcfcf")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV_0\(4),
dataf => \GRLFPC2_0.N_1570\,
datae => \GRLFPC2_0.R.FSR.TEM\(4),
datad => \GRLFPC2_0.R.I.EXC\(4),
datac => \GRLFPC2_0.N_1517\,
datab => N_407);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_0_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfc0c0c0cfcfcfcf")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV_0\(3),
dataf => \GRLFPC2_0.N_1570\,
datae => \GRLFPC2_0.R.FSR.TEM\(3),
datad => \GRLFPC2_0.R.I.EXC\(3),
datac => \GRLFPC2_0.N_1517\,
datab => N_406);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_0_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfc0c0c0cfcfcfcf")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV_0\(2),
dataf => \GRLFPC2_0.N_1570\,
datae => \GRLFPC2_0.R.FSR.TEM\(2),
datad => \GRLFPC2_0.R.I.EXC\(2),
datac => \GRLFPC2_0.N_1517\,
datab => N_405);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_76_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333ffff333fffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7272\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_237\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(61));
\GRLFPC2_0_R_STATE_RNO_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000303030")
port map (
combout => \GRLFPC2_0.R.STATE_0_0_0__G1\,
dataf => \GRLFPC2_0.N_1309\,
datae => CPO_EXCZ,
datad => N_11,
datac => N_7,
datab => \GRLFPC2_0.N_1669\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffff0fff00")
port map (
combout => N_35959,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(21),
datae => \GRLFPC2_0.R.FSR.RD\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(2));
GRLFPC2_0_R_MK_BUSY_RET_4_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000000000000000")
port map (
combout => \GRLFPC2_0.N_2115\,
dataf => \GRLFPC2_0.FPO.BUSY_O\,
datae => \GRLFPC2_0.R.MK.RST_4\,
datad => \GRLFPC2_0.HOLDN_O\,
datac => \GRLFPC2_0.R.MK.HOLDN2_O\,
datab => N_7);
\GRLFPC2_0_V_FSR_FTT_1_IV_I_1_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f3f0f3c0")
port map (
combout => \GRLFPC2_0.N_50_1\,
dataf => \GRLFPC2_0.N_1570\,
datae => \GRLFPC2_0.V.FSR.FTT_1_SQMUXA_1\,
datad => \GRLFPC2_0.R.X.SEQERR\,
datac => \GRLFPC2_0.R.FSR.FTT\(2),
datab => \GRLFPC2_0.N_1105\);
\GRLFPC2_0_R_I_EXC_RNO_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f0000000000000")
port map (
combout => \GRLFPC2_0.R.I.EXC_2_0_2__G2\,
dataf => \GRLFPC2_0.R.I.EXC_MB\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(40),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(38));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_SA_I_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc3f03cffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1_0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_I_7_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfcf0000cfff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_7\(31),
dataf => N_31999_1,
datae => N_31918,
datad => N_32066_2,
datac => N_31769_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_15_0_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff00cf00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_15_0\(31),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_7\(31),
datae => N_32739,
datad => N_32279_3,
datac => N_32070_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_I_21_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3ff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_21\(31),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_15_0\(31),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_9_0\(31),
datad => N_31925_1,
datac => N_32438_1,
datab => N_31813_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_I_6_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff0000fffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_6\(31),
dataf => N_31886_2,
datae => N_31945,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_320\,
datac => N_32632_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_I_5_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000003cffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_5\(31),
dataf => N_31919,
datae => N_31766_2,
datad => N_31924_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_I_12_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000cf000000ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_12\(31),
dataf => N_31919_1,
datae => N_31944,
datad => N_31946,
datac => N_32487_2,
datab => N_31892);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_I_19_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffc0000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_19\(31),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_3\(31),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_12\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_9_TZ\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_320\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_I_23_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_23\(31),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_19\(31),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_5\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_6\(31),
datac => N_31922,
datab => N_31929,
dataa => N_31931);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_I_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"4000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__I0_I_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_23\(31),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_21\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_0\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_10\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_1\(31),
dataa => N_31921);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_8_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_8\(11),
dataf => N_27929_1,
datae => N_32046,
datad => N_32023,
datac => N_31819_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_9_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f3ffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_9\(47),
dataf => N_32621,
datae => N_32487_2,
datad => N_32131_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_6_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffffcfff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_6\(47),
dataf => N_32625,
datae => N_28030_I,
datad => N_28580_1,
datac => N_31723_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_13_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"003f00ff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_13\(47),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_6\(47),
datae => N_32340_1,
datad => N_32994,
datac => N_32124_2,
datab => N_32048_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_12_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f300ff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_12\(47),
dataf => N_52556,
datae => N_32340_1,
datad => N_32626,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_320\,
datab => N_31715_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_22_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_22\(47),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_13\(47),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_12\(47),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_9\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_0\(47),
datab => N_32624,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2302\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_2_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000fcffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_2\(47),
dataf => N_32622,
datae => N_32142_1,
datad => N_32434_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_10_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cf00ff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_10\(47),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_2\(47),
datae => N_32340_1,
datad => N_32641,
datac => N_32632_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_23_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"2000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_23\(47),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_15\(47),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_3\(47),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_4\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_17\(47),
datab => N_32620,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_729\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_48__I0_I_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_22\(47),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_23\(47),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2114\);
GRLFPC2_0_COMB_LOCK_1_0_A2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000300000000")
port map (
combout => CPO_LDLOCKZ,
dataf => \GRLFPC2_0.COMB.LOCKGEN.LOCKI_I_I\,
datae => N_85,
datad => \GRLFPC2_0.R.STATE\(1),
datac => \GRLFPC2_0.R.STATE\(0),
datab => N_84);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_A30_7_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000c000000000")
port map (
combout => N_31926,
dataf => N_32487_2,
datae => N_32775_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_A30_26_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000c")
port map (
combout => N_31945,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_320\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(81),
datad => N_31892,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_A26_23_0_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_A26_23_0\(11),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_A29_6_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00000000000000")
port map (
combout => N_32625,
dataf => N_32343_1,
datae => N_33298,
datad => N_31715_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_A29_9_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => N_32628,
dataf => N_28030_I,
datae => N_31768_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIOCHD_64_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1780_I\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3926\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(68),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(64));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_63_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffc0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1811\,
datae => N_32141_1,
datad => N_31715_1,
datac => N_31924_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_0_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cc00300000000000")
port map (
combout => N_33311,
dataf => N_32141_1_0,
datae => N_33298,
datad => N_31768_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff30000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_2\,
dataf => N_33311,
datae => N_27929_1,
datad => N_32230,
datac => N_32093,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_5_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f00000003000")
port map (
combout => N_33316,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(81),
datae => N_33040,
datad => N_32230,
datac => N_31723_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ffff0300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_1\,
dataf => N_31919_1,
datae => N_33316,
datad => N_31762_1,
datac => N_33040,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_1\,
datac => N_33312,
datab => N_33310,
dataa => N_52547);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_10_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcccf000cccc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_15\,
dataf => N_31725_1,
datae => N_32932,
datad => N_33064_1,
datac => N_32120_1,
datab => N_31941_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_14\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_1\,
datad => N_33072,
datac => N_32645_3,
datab => N_31766_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff030ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_4\,
dataf => N_32141_1,
datae => N_33075,
datad => N_33043_I,
datac => N_33057_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_21\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_12\,
datae => N_33055,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_8\,
datab => N_33144);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_21\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_14\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_20\,
datac => N_33064,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_9\,
dataa => N_33058);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_3_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000003000000")
port map (
combout => N_32275,
dataf => N_31886_2,
datae => N_32124_2,
datad => N_31763_1,
datac => N_31813_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_15_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000000000000000")
port map (
combout => N_32287,
dataf => N_31921_1_0,
datae => N_33063_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_2_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccc0000000000000")
port map (
combout => N_32274,
dataf => N_32141_1_0,
datae => N_32052_1,
datad => N_33063_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_8_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000c0000000000")
port map (
combout => N_32280,
dataf => N_32435_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(81),
datad => N_33071_1,
datac => N_31941_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f333f000f000f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_8\,
dataf => N_31725_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_10_3\(59),
datad => N_32246,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A21_0\(59),
datab => N_32048_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_16\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_11\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_10\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_9\,
datab => N_32277);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff3000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_7\,
dataf => N_31886_2,
datae => N_32691,
datad => N_28580_1,
datac => N_31774_1,
datab => N_31808_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_14\,
dataf => N_32700,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_7\,
datad => N_31921_1,
datac => N_32438_1,
datab => N_31941_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333030333300000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_13\,
dataf => N_32712_3,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_6_1\(58),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O27_1_0_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O27_1_0\(58),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_7_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030300000000000")
port map (
combout => N_32695,
dataf => N_31886_2,
datae => N_32142_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O27_1_0\(58),
datac => N_31808_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffff30ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_12\,
dataf => N_32695,
datae => N_31921_1,
datad => N_32702,
datac => N_32705_1,
datab => N_33298);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff303030ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_2\,
dataf => N_31886_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_15_0\(58),
datad => N_31724_1,
datac => N_32425_1,
datab => N_33176);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_16\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_3\,
datad => N_33145_4,
datac => N_31941_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff8")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_20\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_16\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_12\,
datad => N_32710,
datac => N_32432,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_2_0\(58),
dataa => N_31941_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_1_1_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00003f3000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_1_1\(58),
dataf => N_32425_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff3f0f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_19\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_15\,
datae => N_31921_3,
datad => N_32530_I,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_20\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_19\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_14\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_13\,
datab => N_32688,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2063\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_5_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000300000")
port map (
combout => N_32200,
dataf => N_28030_I,
datae => N_28580_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_4_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c0c0c00000000000")
port map (
combout => N_32199,
dataf => N_33138_1,
datae => N_31766_1,
datad => N_32230,
datac => N_31813_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff8")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_23\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_17\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_16\,
datad => N_32196,
datac => N_33145,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_22_0\(57),
dataa => N_32217_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_19\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_13\,
datad => N_32209,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_6\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_23\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_19\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_4\,
datac => N_32195,
datab => N_32197,
dataa => N_32194);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_9_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_6\,
dataf => N_32424,
datae => N_33138_1,
datad => N_31766_1,
datac => N_31989_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_14\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_6\,
datae => N_32425,
datad => N_31921_1,
datac => N_32066_2,
datab => N_32048_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A28_34_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0f000000000000")
port map (
combout => N_32421,
dataf => N_31865_1,
datae => N_32015_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff30030000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_10\,
dataf => N_32341,
datae => N_32498_4,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_11_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c30000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(81),
datae => N_31763_1,
datad => N_32015_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffc00c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_20\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_10\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_15\,
datad => N_31688,
datac => N_31763_1,
datab => N_32418_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff80")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_24\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_17\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_20\,
datac => N_32344_1,
datab => N_31766_1,
dataa => N_32404);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffc000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_6\,
dataf => N_32739,
datae => N_32770,
datad => N_31940_1,
datac => N_31941_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff30000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_5\,
dataf => N_32777,
datae => N_31839_1,
datad => N_32673_I,
datac => N_31924_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_8_1_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3000000c0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A24_8_1\(55),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(81),
datae => N_33071_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_9_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c3000000000000")
port map (
combout => N_32775,
dataf => N_31921_1_0,
datae => N_32775_1,
datad => N_33298,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_0_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0c0000000000000")
port map (
combout => N_32766,
dataf => N_32708_2,
datae => N_31768_1,
datad => N_31864_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_18\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_9\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_10\,
datad => N_32773,
datac => N_32765,
datab => N_32766,
dataa => N_32775);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_11\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_18\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_17\,
datac => N_32784,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2274\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_30_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c000f0000000000")
port map (
combout => N_32552,
dataf => N_32142_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(81),
datad => N_32220_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_29_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"030c000000000000")
port map (
combout => N_32551,
dataf => N_32272_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(81),
datad => N_32136_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_31_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc00000000000000")
port map (
combout => N_32553,
dataf => N_32142_1,
datae => N_32124_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_26_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0003000000000000")
port map (
combout => N_32548,
dataf => N_31819_1,
datae => N_32136_2,
datad => N_32530_I,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_14\,
dataf => N_32548,
datae => N_32553,
datad => N_32552,
datac => N_32551);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf0cc0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_5\,
dataf => N_31819_1,
datae => N_28580_1,
datad => N_33076_1,
datac => N_31899_I,
datab => N_31924_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_37_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c300000000000000")
port map (
combout => N_32559,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(81),
datae => N_31766_2,
datad => N_31769_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_24_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0c0000000c0000")
port map (
combout => N_32546,
dataf => N_31919_1,
datae => N_31766_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_42_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300000000000000")
port map (
combout => N_32564,
dataf => N_32203_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(81),
datad => N_32015_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff3000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_3\,
dataf => N_31819_1,
datae => N_32564,
datad => N_32203_1,
datac => N_32434_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_17\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_5\,
datac => N_32546,
datab => N_32559);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_23_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000c300000")
port map (
combout => N_32545,
dataf => N_32020,
datae => N_32136_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_44_0_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_44_0\(54),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_36_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0030000000000000")
port map (
combout => N_32558,
dataf => N_33076_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(81),
datad => N_31899_I,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_38_0_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f000f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_38_0\(54),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_25_1_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_25_1\(54),
dataf => N_33076_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_10_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0c0c0c03000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_25_1\(54),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_38_0\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_39_0_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff0000ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_39_0\(54),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_16_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => N_32853,
dataf => N_32438_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(81),
datad => N_32047_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff03000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_5\,
dataf => N_32836,
datae => N_31724_1,
datad => N_31775_1,
datac => N_32908_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcccf000cccc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_4\,
dataf => N_31921_1,
datae => N_33141_2,
datad => N_31724_1,
datac => N_32066_2,
datab => N_32069_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_12_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000c")
port map (
combout => N_32849,
dataf => N_31724_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(81),
datad => N_33176,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_9_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffc0300000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_0\,
dataf => N_32849,
datae => N_27297_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(81),
datac => N_32908_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffc300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_14\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_9\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_3\,
datad => N_32839_3,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffce")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_17\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_14\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_4\,
datad => N_32846,
datac => N_31921_1,
datab => N_32838,
dataa => N_32840_3);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff80")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_17\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_13\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_12\,
datac => N_31766_1,
datab => N_31996_1,
dataa => N_32418_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_5_2_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f000000fff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_5_2\(52),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_3_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cc0f000000000000")
port map (
combout => N_33130,
dataf => N_32343_1,
datae => N_32050_1,
datad => N_31765_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_10_0\,
dataf => N_33131,
datae => N_33130,
datad => N_33129,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_22_1\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_22_0\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff30c00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_2\,
dataf => N_33136,
datae => N_33141_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffc0c30000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_9\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_12_TZ\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_13_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c00000000000000")
port map (
combout => N_33140,
dataf => N_31886_2,
datae => N_32705_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_7_0_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3033033300000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_7_0\(52),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_9\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_14\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_10_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_16\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_13\,
dataa => N_33145);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_10\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_255\,
datac => N_32134_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00c000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_4\,
dataf => N_32141_1,
datae => N_33271,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_320\,
datac => N_32120_1,
datab => N_32394_I);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_12\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_13\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_10\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_11\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_9\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2367\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_9_0_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_9_0\(50),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffcc00fffffcf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_255\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2354\,
datad => N_32217_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2767\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2693\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffcf0cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_9\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8695\,
datae => N_32925_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2763\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2505\,
datab => N_31924_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_11_0_49_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff0000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_11_0\(49),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffcf0cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2354\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2648\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_11_0\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_11_1\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2636\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff0c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_13\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1937\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2373\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(81),
datab => N_33206);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffc0c0c0ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_1\,
dataf => N_31725_1,
datae => N_31925_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2499\,
datac => N_33064_1,
datab => N_32120_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff3c000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_1\,
datae => N_32344_1,
datad => N_33063_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_12\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9079\,
datad => N_32344_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2634\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2659\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff0c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_11\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2321\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_255\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2657\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffa8")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_12\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_13\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_11\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2725\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2602\,
dataa => N_31763_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_35_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300000000000000")
port map (
combout => N_32357,
dataf => N_32550_1,
datae => N_32632_1,
datad => N_32124_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_32_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000003300000")
port map (
combout => N_32354,
dataf => N_33040,
datae => N_32015_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_49_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff3003ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_31_1\(48),
datae => N_32354,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_19_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000c00000000000")
port map (
combout => N_32341,
dataf => N_31940_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(81),
datad => N_31989_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83),
datab => N_32140_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_49_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_5\,
dataf => N_32340,
datae => N_32343,
datad => N_32341);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_26_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f30000000f000000")
port map (
combout => N_32348,
dataf => N_33136_1,
datae => N_32632_1,
datad => N_32705_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_24_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000303f00000000")
port map (
combout => N_32346,
dataf => N_32925_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_247\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_23_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03cf000000000000")
port map (
combout => N_32345,
dataf => N_32345_2,
datae => N_33057_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_49_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_12\,
dataf => N_32346,
datae => N_32345,
datad => N_32336,
datac => N_32272_2,
datab => N_31765_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_49_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_15\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_12\,
datae => N_33136_1,
datad => N_31766_1,
datac => N_32418_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_49_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_15\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_7\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_13\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_6\,
dataa => N_33067);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_45_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_354\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2648\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2622_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_44_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffcf0cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_44__G2_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2263\,
datae => N_31921_3,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2703\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2498\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2508\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_3_0_41_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3_0\(41),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_40_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_40__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_450\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_523\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_1_0\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1932\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2572\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_39_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_39__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1042\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_450\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_39__G2_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_1_0\(39),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2572\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_37_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffc0c0ffffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_450\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_346\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2300\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2658\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_38_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffcf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_450\,
datae => N_31725_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2490\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2518\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2546\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_38_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2_3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1042\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2689\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2505\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3f0f33000f0f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_4\,
dataf => N_31725_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2526\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2508\,
datac => N_32645_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_10\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8752\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_4\,
datad => N_31725_1,
datac => N_32203_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2525\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_14\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_10\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2114\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2703\,
datac => N_31763_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2337\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2341\,
datad => N_31921_1,
datac => N_31811_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffff0f03000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_16\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_13\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2671\,
datad => N_33143_1,
datac => N_32438_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff2")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_16\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_14\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_445\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2706\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_35_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffcf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_35__G2_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2405\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2300\,
datad => N_33001_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2407\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2633\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_35_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_35__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_35__G2_3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_35__G2_2\,
datad => N_32141_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2505\,
datab => N_32048_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_1_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff000000c0000000")
port map (
combout => N_31989,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(81),
datae => N_32069_2,
datad => N_31989_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff8")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_9\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_7\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_8\,
datab => N_33001_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0_0\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff3000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_13\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_0\,
datae => N_33274,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datac => N_32418_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A24_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000c000c0000000")
port map (
combout => N_33255,
dataf => N_32289_2,
datae => N_32064_1,
datad => N_31723_1,
datac => N_32220_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_12\,
dataf => N_33276,
datae => N_33255,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_9_0\(62),
datac => N_33136_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_15\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_13\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_14\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_16\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_12\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2586\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_21_RNI4CMFC_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffc0ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_7\,
dataf => N_32487,
datae => N_31921_1,
datad => N_32497,
datac => N_32500_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_26_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000003c00000000")
port map (
combout => N_32492,
dataf => N_31921_1_0,
datae => N_33232,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_26_RNI2OHE9_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffc3ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_10\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_6_TZ\,
datad => N_32492,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_30_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => N_32496,
dataf => N_32775_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(81),
datad => N_32015_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_18_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0033003000000000")
port map (
combout => N_32484,
dataf => N_32141_1_0,
datae => N_32775_1,
datad => N_33232,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A20_RNIM89BH1_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_10\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_8\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_7\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_4\,
datab => N_32483,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_5_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_30_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c0000c00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2419\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2526\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf0f0f0cc000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2_1\,
dataf => N_32619_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2485\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2536\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2546\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffc0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2_1\,
datae => N_27776_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datac => N_32069_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1931\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2283\,
datad => N_32020,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2485\,
datab => N_32885_I);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff3000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_3\,
dataf => N_31768,
datae => N_31769,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A9_0_1\(28),
datac => N_31763_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A9_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03cc000000030000")
port map (
combout => N_31762,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2_1\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffc00000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_2\,
dataf => N_31762,
datae => N_32131_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datac => N_31766_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A9_3_0\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_4_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c300000000000000")
port map (
combout => N_31767,
dataf => N_31819_1,
datae => N_31763_1,
datad => N_31767_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00c00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_1\,
dataf => N_31767,
datae => N_32032_I,
datad => N_32142_1,
datac => N_31765_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff80")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_2\,
datac => N_31925_1,
datab => N_32131_1,
dataa => N_31753);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_11_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3003000000000000")
port map (
combout => N_32912,
dataf => N_32070_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_13_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c300000000000000")
port map (
combout => N_32914,
dataf => N_32620_1,
datae => N_28580_1,
datad => N_32050_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_4_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0cf000000000000")
port map (
combout => N_32905,
dataf => N_32708_2,
datae => N_32220_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_12_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"003c000000000000")
port map (
combout => N_32913,
dataf => N_31921_1_0,
datae => N_31766_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_13_0\,
dataf => N_32905,
datae => N_32913,
datad => N_32908,
datac => N_32932,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_13_TZ\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcccf000cccc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_6\,
dataf => N_31921_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_1_TZ\,
datad => N_31766_1,
datac => N_31838_1,
datab => N_31941_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_20\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_13_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_6\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_11\,
dataa => N_32904);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffff3f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_9\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8752\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2796\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_10_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000030000000000")
port map (
combout => N_31819,
dataf => N_31819_1,
datae => N_31899_I,
datad => N_31819_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_4_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c3000000000000")
port map (
combout => N_31813,
dataf => N_31725_1_0,
datae => N_31813_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_3\,
dataf => N_31819,
datae => N_31813,
datad => N_31817,
datac => N_31814);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffff0003000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_5\,
dataf => N_31810,
datae => N_33138_1,
datad => N_31811_2,
datac => N_32136_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_5\,
datac => N_31808,
datab => N_31809,
dataa => N_31818);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_24_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffc000c000c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_24__G2_0\,
dataf => N_33069,
datae => N_32487_2,
datad => N_31762_1,
datac => N_31808_1,
datab => N_33023);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_21_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffcccf000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_21__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1922\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2779\,
datad => N_32344_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2551\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_7_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000030000")
port map (
combout => N_32127,
dataf => N_31921_1_0,
datae => N_31768_1,
datad => N_33040,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_7_RNIGSG04_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff03000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_7\,
dataf => N_32127,
datae => N_27929_1,
datad => N_32093,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_2_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03cf000000000000")
port map (
combout => N_32122,
dataf => N_32620_1,
datae => N_31769_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_0_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c33000000000000")
port map (
combout => N_32120,
dataf => N_32620_1,
datae => N_32120_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_13_RNIJ16K5_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_15_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_2\,
datae => N_32133,
datad => N_32143,
datac => N_32124,
datab => N_32141);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_9_0_RNIQL7JK1_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff8")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_17\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_15_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_11\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_14\,
datab => N_31921_3,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_9_0\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_4_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000300000000")
port map (
combout => N_31867,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(81),
datae => N_33298,
datad => N_31819_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_3_0_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f0f0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_3_0\(18),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A15_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c0c0c000c0c00000")
port map (
combout => N_31862,
dataf => N_31886_2,
datae => N_31887,
datad => N_28580_1,
datac => N_31774_1,
datab => N_31808_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_9\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_2_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_3\,
datac => N_31862,
datab => N_31875,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_9_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000c00000000000")
port map (
combout => N_31719,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(81),
datae => N_32673_I,
datad => N_33136_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_9_RNISC2D2_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffc000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_0\,
dataf => N_31886_2,
datae => N_31719,
datad => N_32566_1,
datac => N_31691_I,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O18_2_RNIQ0TD3_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00000300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_3\,
dataf => N_31709,
datae => N_31688,
datad => N_31703,
datac => N_33176,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_6_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000c0000000")
port map (
combout => N_31716,
dataf => N_31921_1_0,
datae => N_32069_2,
datad => N_33136_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_4_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000003c0000")
port map (
combout => N_31714,
dataf => N_31688,
datae => N_32688_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_2_0_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_2_0\(17),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_2_0_RNIHO1C3_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00f00030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_1_0\,
dataf => N_31714,
datae => N_32550_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_247\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_2_0\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O18_3_RNIVC6U7_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_1_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_2\,
datad => N_31713,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_0_0\(17),
datab => N_31704);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_8\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_9\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1937\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2581\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2063\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1941\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_O2_RNI6STA4_39_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_16__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_523\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_16__G2_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_16__G2_1\,
datac => N_32925_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2505\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_14_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffcfff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_14__G2\,
dataf => N_33148,
datae => N_33133_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2214\,
datac => N_52211,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2659\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_2_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00003c0000000000")
port map (
combout => N_33198,
dataf => N_32632_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(81),
datad => N_32705_1,
datac => N_33176,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_4_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c0000c0000000000")
port map (
combout => N_33200,
dataf => N_32708_2,
datae => N_32632_1,
datad => N_31864_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_13_RNIPQNS_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_7\,
dataf => N_33200,
datae => N_33202,
datad => N_33203,
datac => N_33198,
datab => N_33209);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_35_RNIPMMN3_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffc0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2063\,
datae => N_27776_2,
datad => N_32069_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_8__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_8__G2_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1941\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2359\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1967_1\,
datab => N_32136_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cc000000fcf0f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_255\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2490\,
datad => N_31762_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_15_0\(7),
datab => N_31808_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_8\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_726\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2288\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2290\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_7_1_0_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0cc00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_7_1\(6),
dataf => N_32052_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffccc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_12\,
dataf => N_32985,
datae => N_32980,
datad => N_32995_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_8_0\(6),
datab => N_33023);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffc0ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_11\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_4\,
datae => N_31921_1,
datad => N_32991,
datac => N_32203_1,
datab => N_31813_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_17\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_12\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_7\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2373\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_11\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2268\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_6\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2267\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_5\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2581\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A3_RNIM9H52_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8994\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1982\,
datad => N_32662_I,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2636\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_1_RNIV2205_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_10\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_4\,
datad => N_33001_1,
datac => N_31838_1,
datab => N_31924_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_13_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000300000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1958\,
dataf => N_31921_1_0,
datae => N_31996_1,
datad => N_32136_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_RNI3BIAP_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_11\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_10\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1937\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_13\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1954\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_21_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => N_33148,
dataf => N_32438_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(81),
datad => N_32688_1,
datac => N_32047_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_0_0_RNI3RJD_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcccf000cccc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2_1\,
dataf => N_33133_1,
datae => N_32128_1,
datad => N_31763_1,
datac => N_31762_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_0_RNI4RIS5_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8639\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9471\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_596\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_2__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19\(9),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2214\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2598\,
datac => N_27776_2,
datab => N_31941_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000c000ffffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_1__G2_0\,
dataf => N_31919_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2784\,
datad => N_27776_2,
datac => N_32069_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_1__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8639\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_1__G2_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1941\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1940\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_6_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000000000000000")
port map (
combout => N_33359,
dataf => N_32340_1_0,
datae => N_31941_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_3_RNICLS43_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_3\,
dataf => N_33359,
datae => N_33356,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A12_0_0\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_247\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82));
GRLFPC2_0_R_A_LD_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000cf000000")
port map (
combout => \GRLFPC2_0.R.A.LD_0_0_G1\,
dataf => \GRLFPC2_0.COMB.LOCKGEN.LOCKI_I_I\,
datae => \GRLFPC2_0.N_939_I_0_A2_2\,
datad => \GRLFPC2_0.R.A.LD_0_0_G1_0\,
datac => N_70,
datab => N_69);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A3_6_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f000003000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2474\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2457\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_377\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(73),
datab => N_56);
\GRLFPC2_0_R_A_RF1REN_RNO_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300000000000000")
port map (
combout => N_36379,
dataf => \GRLFPC2_0.COMB.LOCKGEN.LOCKI_I_1\,
datae => \GRLFPC2_0.COMB.V.A.RF1REN_1_0_7636_I_1\,
datad => N_73,
datac => N_72,
datab => N_36289);
GRLFPC2_0_COMB_UN6_IUEXEC_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f3000000ff0000")
port map (
combout => \GRLFPC2_0.COMB.UN6_IUEXEC_1\,
dataf => \GRLFPC2_0.R.MK.BUSY_4\,
datae => \GRLFPC2_0.R.MK.BUSY_O\,
datad => \GRLFPC2_0.COMB.ANNULFPU_1_O_0\,
datac => \GRLFPC2_0.R.MK.RST_O_0\,
datab => \GRLFPC2_0.R.MK.HOLDN2_O_0\);
GRLFPC2_0_COMB_UN6_IUEXEC: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f00000000")
port map (
combout => \GRLFPC2_0.N_1255\,
dataf => \GRLFPC2_0.COMB.UN6_IUEXEC_1\,
datae => \GRLFPC2_0.R.MK.RST\,
datad => \GRLFPC2_0.N_178\,
datac => \GRLFPC2_0.R.MK.RST2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_15_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000c000")
port map (
combout => N_32852,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_320\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(81),
datad => N_32908_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_11_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000c00000000000")
port map (
combout => N_32848,
dataf => N_32066_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(81),
datad => N_33176,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_5_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c0c0c00000000000")
port map (
combout => N_32693,
dataf => N_31839_1,
datae => N_32064_1,
datad => N_32566_1,
datac => N_31767_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_2_0_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0030333000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_2_0\(58),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_A30_0_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc000c0000000000")
port map (
combout => N_31919,
dataf => N_31919_1,
datae => N_31892,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(78));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_OPREXCSHFT_UN14_EXMIPTRLSBS_RNI0FGR1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000c00000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3729_I_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5065\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN14_EXMIPTRLSBS\);
\GRLFPC2_0_R_A_RF1REN_RNO_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f000ff00")
port map (
combout => N_36380,
dataf => \GRLFPC2_0.COMB.LOCKGEN.LOCKI_I_I\,
datae => N_36304,
datad => \GRLFPC2_0.COMB.RS1V_1\,
datac => \GRLFPC2_0.COMB.RS1D_1\);
\GRLFPC2_0_R_A_RF2REN_RNO_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff00f000")
port map (
combout => N_36382,
dataf => \GRLFPC2_0.COMB.LOCKGEN.LOCKI_I_I\,
datae => N_36304,
datad => \GRLFPC2_0.COMB.RS1V_1\,
datac => \GRLFPC2_0.COMB.RS1D_1\);
\GRLFPC2_0_R_I_EXC_RNO_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000003000")
port map (
combout => \GRLFPC2_0.R.I.EXC_2_0_1__G2\,
dataf => \GRLFPC2_0.N_1470\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(40),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(38),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(41));
\GRLFPC2_0_R_I_EXC_RNO_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000f0")
port map (
combout => \GRLFPC2_0.R.I.EXC_2_0_3__G2\,
dataf => \GRLFPC2_0.N_1470\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(40),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(38));
\GRLFPC2_0_R_I_EXC_RNO_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000cc00c000")
port map (
combout => \GRLFPC2_0.R.I.EXC_2_0_4__G2\,
dataf => \GRLFPC2_0.N_1470\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(40),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(38),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(41));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_40_RNIKSJ6C: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc0000cc0f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_1_TZ\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
GRLFPC2_0_R_X_FPOP_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000000")
port map (
combout => \GRLFPC2_0.R.X.FPOP_0_0_G1\,
dataf => \GRLFPC2_0.R.M.FPOP\,
datae => N_291,
datad => N_292);
GRLFPC2_0_R_X_LD_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000000")
port map (
combout => \GRLFPC2_0.R.X.LD_0_0_G1\,
dataf => \GRLFPC2_0.R.M.LD\,
datae => N_291,
datad => N_292);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7260\,
dataf => N_57,
datae => N_61,
datad => N_59,
datac => N_62);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7259\,
dataf => N_57,
datae => N_61,
datad => N_59,
datac => N_62);
GRLFPC2_0_R_M_AFQ_RET_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.R.M.AFQ_RET_0_0_G1\,
dataf => \GRLFPC2_0.N_1830_O\,
datae => \GRLFPC2_0.R.A.AFQ_O\);
GRLFPC2_0_R_M_AFSR_RET_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.R.M.AFSR_RET_0_0_G1\,
dataf => \GRLFPC2_0.N_1830_O\,
datae => \GRLFPC2_0.R.A.AFSR_O\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4459\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_RNIDSCN5_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f000f0f0f000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(58),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(58),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_317__G1\,
datac => \GRLFPC2_0.FPI.LDOP_4\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0ff0f000ffff00")
port map (
combout => N_58821,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_58820,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(310));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0ff0f000ffff00")
port map (
combout => N_58746,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_9_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_58745,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(306));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0ff0f000ffff00")
port map (
combout => N_58723,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_58722,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(307));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0ff0f000ffff00")
port map (
combout => N_58700,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_58699,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(308));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0ff0f000ffff00")
port map (
combout => N_58677,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_58676,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(309));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0f0ff0f00ff0f0")
port map (
combout => N_58657,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff0ff0ff000ff0")
port map (
combout => N_58632,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_58631,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(259));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ffff000f0ff0f0")
port map (
combout => N_58609,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_58608,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(260));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0ff0f000ffff00")
port map (
combout => N_58586,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_58585,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(261));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff0ff0ff000ff0")
port map (
combout => N_58561,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_24_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_58560,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(291));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff000ff0ff0ff00")
port map (
combout => N_58538,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_23_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_58537,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(292));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0ff00f0ff0f0f0")
port map (
combout => N_58515,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_22_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_58514,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(293));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff0ff0ff000ff0")
port map (
combout => N_58492,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_21_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_58491,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(294));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff000ff0ff0ff00")
port map (
combout => N_58469,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_20_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_58468,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(295));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0ff00f0ff0f0f0")
port map (
combout => N_58446,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_58445,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(296));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0f0ff0f00ff0f0")
port map (
combout => N_58423,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_58422,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(297));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0f0ff0f0f00ff0")
port map (
combout => N_58400,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_58399,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(298));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff00ff00f0ff0f0")
port map (
combout => N_58377,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_16_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_58376,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(299));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ffff000ff00ff0")
port map (
combout => N_58354,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_15_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_58353,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(300));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff00ff000ffff00")
port map (
combout => N_58331,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_14_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_58330,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(301));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0ff0f00ff00ff0")
port map (
combout => N_58308,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_58307,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(302));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff00ff00f0ff0f0")
port map (
combout => N_58285,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_12_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_58284,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(303));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff00ff00f0ff0f0")
port map (
combout => N_58262,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_58261,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(304));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ffff000ff00ff0")
port map (
combout => N_58239,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_10_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_58238,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(305));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ffff000ff00ff0")
port map (
combout => N_58216,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_39_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_58215,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(276));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0ff0f000ffff00")
port map (
combout => N_58193,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_38_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_58192,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(277));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff00ff000ffff00")
port map (
combout => N_58170,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_37_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_58169,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(278));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff00ff00f0ff0f0")
port map (
combout => N_58147,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_58146,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(279));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ffff000ff00ff0")
port map (
combout => N_58124,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_35_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_58123,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(280));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0ff0f000ffff00")
port map (
combout => N_58101,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_58100,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(281));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff00ff000ffff00")
port map (
combout => N_58078,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_58077,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(282));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff00ff00f0ff0f0")
port map (
combout => N_58055,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_58054,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(283));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff00ff00f0ff0f0")
port map (
combout => N_58032,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_58031,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(284));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff00f0f0ff0f0f0")
port map (
combout => N_58009,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_30_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_58008,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(285));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0ff00f0ff0f0f0")
port map (
combout => N_57986,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_57985,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(286));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0ff00f0ff0f0f0")
port map (
combout => N_57963,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_57962,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(287));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0ff00f0ff0f0f0")
port map (
combout => N_57940,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_57939,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(288));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0ff00f0ff0f0f0")
port map (
combout => N_57917,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_57916,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(289));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0ff00f0ff0f0f0")
port map (
combout => N_57894,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_57893,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(290));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0ff0f000ffff00")
port map (
combout => N_57871,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_57870,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(262));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0ff0f000ffff00")
port map (
combout => N_57848,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_57847,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(263));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ffff000f0ff0f0")
port map (
combout => N_57825,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_57824,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(264));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ffff000f0ff0f0")
port map (
combout => N_57802,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_57801,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(265));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff000ff0ff0ff00")
port map (
combout => N_57779,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_49_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_57778,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(266));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff0ff0ff000ff0")
port map (
combout => N_57756,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_57755,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(267));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0ff0f000ffff00")
port map (
combout => N_57733,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_57732,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(268));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0ff0f000ffff00")
port map (
combout => N_57710,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_46_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_57709,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(269));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff000ff0ff0ff00")
port map (
combout => N_57687,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_45_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_57686,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(270));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff0ff0ff000ff0")
port map (
combout => N_57664,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_44_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_57663,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(271));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff000ff0ff0ff00")
port map (
combout => N_57641,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_43_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_57640,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(272));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff0ff0ff000ff0")
port map (
combout => N_57618,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_42_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_57617,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(273));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff000ff0ff0ff00")
port map (
combout => N_57595,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_41_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_57594,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(274));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0f0ff0f0f00ff0")
port map (
combout => N_57572,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_40_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_57571,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(275));
\GRLFPC2_0_R_A_RF2REN_RNO_0_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000003f003f003f")
port map (
combout => N_36334,
dataf => \GRLFPC2_0.N_889\,
datae => N_50,
datad => \GRLFPC2_0.N_896\,
datac => \GRLFPC2_0.COMB.FPDECODE.RS1D5\,
datab => \GRLFPC2_0.N_884\);
\GRLFPC2_0_R_A_RF1REN_RNO_1_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000fff00000000")
port map (
combout => N_36289,
dataf => N_50,
datae => \GRLFPC2_0.N_896\,
datad => \GRLFPC2_0.COMB.FPDECODE.RS1D5\,
datac => \GRLFPC2_0.N_884\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A12_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3330303000000000")
port map (
combout => N_33352,
dataf => N_32645_3,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_247\,
datad => N_31766_2,
datac => N_33367,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_A30_27_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000c00000000000")
port map (
combout => N_31946,
dataf => N_32066_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(81),
datad => N_32015_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_233_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cf000000c000")
port map (
combout => N_36374,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\(11),
datae => \GRLFPC2_0.FPI.LDOP_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7612_I_1_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIHKHD_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7612_I_1_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
datae => \GRLFPC2_0.R.MK.RST2\,
datad => N_7);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_232_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cf000000c000")
port map (
combout => N_36375,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\(12),
datae => \GRLFPC2_0.FPI.LDOP_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7612_I_1_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(245));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c0ff0000c03000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_13_TZ\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_9_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cf0fc000c000c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_1_TZ\,
dataf => N_27297_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datad => N_32272_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_4_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fff0fcfffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_I_0_4\(11),
dataf => N_27929_1,
datae => N_33298,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A28_24_0\(60),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_I_9_TZ_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0fffffffff0ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_9_TZ\(31),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_12_RNO_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccfffcffcfffffff")
port map (
combout => N_52556,
dataf => N_31999_1,
datae => N_32708_2,
datad => N_32120_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000003c0000000")
port map (
combout => N_52547_TZ,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_316_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffccc0fcc0fccc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_316__G1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1281_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_58\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7035\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7051\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_3_RNISFVF5: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffccc0fcc0fccc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_317__G1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1281_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_58\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7035\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7034\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_CIN_3_RNI3MFN3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffccc0fcc0fccc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_318__G1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1281_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_58\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN_3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN12_SRTOSTICKY_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN12_SRTOSTICKY_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(9),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_O3_2_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0fff0f0cffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN11_WQSTSETS\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_112_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(112),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datae => N_663);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_111_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(111),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datae => N_664);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_110_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(110),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datae => N_665);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_109_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(109),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datae => N_666);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_108_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(108),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datae => N_667);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_107_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(107),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datae => N_668);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_106_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(106),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datae => N_669);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_105_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(105),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datae => N_670);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_104_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(104),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datae => N_671);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_103_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(103),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datae => N_672);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_102_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(102),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datae => N_673);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_101_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(101),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datae => N_674);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_100_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(100),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datae => N_675);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_99_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(99),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datae => N_676);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_98_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(98),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datae => N_677);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_97_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(97),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datae => N_678);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_96_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(96),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datae => N_679);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_95_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(95),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datae => N_680);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_94_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(94),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datae => N_681);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_93_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(93),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datae => N_682);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_92_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(92),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datae => N_683);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_91_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(91),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datae => N_684);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_90_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(90),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datae => N_685);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_89_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(89),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datae => N_686);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_88_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(88),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datae => N_687);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_87_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(87),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datae => N_688);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_86_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(86),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datae => N_689);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_85_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(85),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datae => N_690);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_84_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(84),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datae => N_691);
\GRLFPC2_0_R_I_EXC_0_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000048c00008c8c")
port map (
combout => \GRLFPC2_0.R.I.EXC_MB\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_28\,
datae => \GRLFPC2_0.N_1470\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_27\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4664\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4662\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\);
GRLFPC2_0_COMB_V_E_STDATA2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA2\,
dataf => N_151,
datae => N_152);
GRLFPC2_0_COMB_V_A_SEQERR_1_0_A2_0_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000c000000000")
port map (
combout => \GRLFPC2_0.COMB.V.A.SEQERR_1_0_A2_0_3\,
dataf => \GRLFPC2_0.FPCI_O\(62),
datae => \GRLFPC2_0.FPCI_O\(69),
datad => \GRLFPC2_0.FPCI_O\(59),
datac => \GRLFPC2_0.FPCI_O\(60),
datab => \GRLFPC2_0.N_1837_O\);
GRLFPC2_0_COMB_V_A_SEQERR_1_0_O2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0c0c0cff000000")
port map (
combout => \GRLFPC2_0.N_11\,
dataf => \GRLFPC2_0.N_10\,
datae => \GRLFPC2_0.COMB.V.A.SEQERR_1_0_A2_0_3\,
datad => \GRLFPC2_0.N_7\,
datac => \GRLFPC2_0.FPCI_O\(62),
datab => \GRLFPC2_0.FPCI_O\(69));
GRLFPC2_0_WRADDR_0_SQMUXA_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000000000000")
port map (
combout => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
dataf => N_395,
datae => N_396,
datad => N_397);
\GRLFPC2_0_COMB_DBGDATA_4_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffff00f0f0")
port map (
combout => CPO_DBG_DATAZ(17),
dataf => N_397,
datae => N_398,
datad => N_680,
datac => N_616);
\GRLFPC2_0_COMB_DBGDATA_4_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffff00f0f0")
port map (
combout => CPO_DBG_DATAZ(18),
dataf => N_397,
datae => N_398,
datad => N_681,
datac => N_617);
\GRLFPC2_0_COMB_DBGDATA_4_12_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff00f0f0")
port map (
combout => CPO_DBG_DATAZ(12),
dataf => N_397,
datae => N_398,
datad => N_675,
datac => N_611);
\GRLFPC2_0_COMB_DBGDATA_4_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff00f0f0")
port map (
combout => CPO_DBG_DATAZ(28),
dataf => N_397,
datae => N_398,
datad => N_691,
datac => N_627);
\GRLFPC2_0_COMB_V_E_STDATA_1_1_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff00fffff0f0")
port map (
combout => \GRLFPC2_0.N_3156\,
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.R.A.AFSR\,
datad => N_681,
datac => N_617);
\GRLFPC2_0_COMB_DBGDATA_4_15_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff00f0f0")
port map (
combout => CPO_DBG_DATAZ(15),
dataf => N_397,
datae => N_398,
datad => N_678,
datac => N_614);
\GRLFPC2_0_COMB_DBGDATA_4_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff00f0f0")
port map (
combout => CPO_DBG_DATAZ(19),
dataf => N_397,
datae => N_398,
datad => N_682,
datac => N_618);
\GRLFPC2_0_COMB_DBGDATA_4_20_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff00f0f0")
port map (
combout => CPO_DBG_DATAZ(20),
dataf => N_397,
datae => N_398,
datad => N_683,
datac => N_619);
\GRLFPC2_0_COMB_DBGDATA_4_21_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff00f0f0")
port map (
combout => CPO_DBG_DATAZ(21),
dataf => N_397,
datae => N_398,
datad => N_684,
datac => N_620);
\GRLFPC2_0_COMB_DBGDATA_4_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff00f0f0")
port map (
combout => CPO_DBG_DATAZ(29),
dataf => N_397,
datae => N_398,
datad => N_692,
datac => N_628);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNI0DHE1_71_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcfffcfffcfff0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(71));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_258_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0cf3fffff30c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_258__N_5_I\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8_0\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6961\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58));
GRLFPC2_0_COMB_UN1_MEXC_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f00ff0f0fffff")
port map (
combout => \GRLFPC2_0.COMB.UN1_MEXC_1_0\,
dataf => \GRLFPC2_0.R.FSR.TEM\(2),
datae => \GRLFPC2_0.R.FSR.TEM\(3),
datad => \GRLFPC2_0.R.I.EXC\(2),
datac => \GRLFPC2_0.R.I.EXC\(3));
GRLFPC2_0_COMB_UN1_MEXC_1_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f00ff0f0fffff")
port map (
combout => \GRLFPC2_0.COMB.UN1_MEXC_1_1\,
dataf => \GRLFPC2_0.R.FSR.TEM\(0),
datae => \GRLFPC2_0.R.FSR.TEM\(1),
datad => \GRLFPC2_0.R.I.EXC\(0),
datac => \GRLFPC2_0.R.I.EXC\(1));
GRLFPC2_0_COMB_UN1_MEXC_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fff000000000000")
port map (
combout => \GRLFPC2_0.N_1768\,
dataf => \GRLFPC2_0.COMB.UN1_MEXC_1_1\,
datae => \GRLFPC2_0.COMB.UN1_MEXC_1_0\,
datad => \GRLFPC2_0.R.FSR.TEM\(4),
datac => \GRLFPC2_0.R.I.EXC\(4));
\GRLFPC2_0_R_FSR_FTT_RNO_0_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000c0000000c000")
port map (
combout => \GRLFPC2_0.R.FSR.FTT_M_2\(0),
dataf => \GRLFPC2_0.N_1768\,
datae => \GRLFPC2_0.V.FSR.FTT_3_SQMUXA_I_A3_0\,
datad => \GRLFPC2_0.N_3422\,
datac => \GRLFPC2_0.R.FSR.FTT\(0),
datab => N_7);
\GRLFPC2_0_R_FSR_FTT_RNO_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcf0f0ffcc0000")
port map (
combout => \GRLFPC2_0.R.FSR.FTT_0_0_0__G1\,
dataf => \GRLFPC2_0.N_1570\,
datae => \GRLFPC2_0.R.FSR.FTT_M_2\(0),
datad => \GRLFPC2_0.V.FSR.FTT_1_SQMUXA_1\,
datac => N_7,
datab => \GRLFPC2_0.N_1105\);
GRLFPC2_0_R_I_PC_RET_60_RNI7KV4: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => N_9);
\GRLFPC2_0_R_I_RES_RNO_63_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0303ff000c0cff00")
port map (
combout => \GRLFPC2_0.COMB.V.I.RES_1\(63),
dataf => \GRLFPC2_0.FPI.OP2\(63),
datae => \GRLFPC2_0.N_1470\,
datad => \GRLFPC2_0.FPO.SIGN\,
datac => N_127,
datab => N_126);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bcb0bf838c808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10074\,
dataf => \GRLFPC2_0.FPO.FRAC\(49),
datae => \GRLFPC2_0.FPO.FRAC\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_CIN_3_RNI3MFN3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cc333cc33cc333cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1281_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_58\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN_3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bf838cb0bc808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10080\,
dataf => \GRLFPC2_0.FPO.FRAC\(54),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_176__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_15_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bcb0bf838c808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10067\,
dataf => \GRLFPC2_0.FPO.FRAC\(42),
datae => \GRLFPC2_0.FPO.FRAC\(41),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_4_0_RNIJIFB1_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30cf3fc000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7051\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6961\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bcb0bf838c808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10082\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_175__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_257_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfffcf00c0ffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10525\,
dataf => \GRLFPC2_0.FPO.EXP\(1),
datae => \GRLFPC2_0.FPO.EXP\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_254_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10514\,
dataf => \GRLFPC2_0.FPO.EXP\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(241));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_253_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfffcf00c0ffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10529\,
dataf => \GRLFPC2_0.FPO.EXP\(5),
datae => \GRLFPC2_0.FPO.EXP\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(240));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_249_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfffcf00c0ffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10533\,
dataf => \GRLFPC2_0.FPO.EXP\(9),
datae => \GRLFPC2_0.FPO.EXP\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_248_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10520\,
dataf => \GRLFPC2_0.FPO.EXP\(10),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0fff000f0fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_46_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10036\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(46),
datae => \GRLFPC2_0.FPO.FRAC\(11),
datad => \GRLFPC2_0.FPO.FRAC\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M2_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M2\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M12_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0f03ffff0f00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M2\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M12_RNIUT1C_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0f0f00000f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M13\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM12\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc30fc30fc30cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10935\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10939\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcf0fcff0c000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10944\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(241));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bf838cb0bc808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10056\,
dataf => \GRLFPC2_0.FPO.FRAC\(30),
datae => \GRLFPC2_0.FPO.FRAC\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bcb0bf838c808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10076\,
dataf => \GRLFPC2_0.FPO.FRAC\(51),
datae => \GRLFPC2_0.FPO.FRAC\(50),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bf838cb0bc808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075\,
dataf => \GRLFPC2_0.FPO.FRAC\(49),
datae => \GRLFPC2_0.FPO.FRAC\(50),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10014\,
dataf => \GRLFPC2_0.FPI.LDOP_5\,
datae => \GRLFPC2_0.FPI.OP2\(49),
datad => \GRLFPC2_0.FPI.OP2\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(124));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10134\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10014\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_10_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10012\,
dataf => \GRLFPC2_0.FPI.LDOP_5\,
datae => \GRLFPC2_0.FPI.OP2\(47),
datad => \GRLFPC2_0.FPI.OP2\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(126));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_10_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10132\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(10),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10012\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bf838cb0bc808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10055\,
dataf => \GRLFPC2_0.FPO.FRAC\(29),
datae => \GRLFPC2_0.FPO.FRAC\(30),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_23_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bf838cb0bc808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10059\,
dataf => \GRLFPC2_0.FPO.FRAC\(33),
datae => \GRLFPC2_0.FPO.FRAC\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_44_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10038\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(44),
datae => \GRLFPC2_0.FPO.FRAC\(13),
datad => \GRLFPC2_0.FPO.FRAC\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_42_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10040\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(42),
datae => \GRLFPC2_0.FPO.FRAC\(15),
datad => \GRLFPC2_0.FPO.FRAC\(14),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_43_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10039\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(43),
datae => \GRLFPC2_0.FPO.FRAC\(14),
datad => \GRLFPC2_0.FPO.FRAC\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_45_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9977\,
dataf => \GRLFPC2_0.FPI.LDOP_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(161),
datac => N_704);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_45_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10097\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(45),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9977\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_45_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3ff333fc0cc000c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(45),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(12),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(46),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_46_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9976\,
dataf => \GRLFPC2_0.FPI.LDOP_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(162),
datac => N_703);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_46_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10096\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(46),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9976\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_46_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3ff333cc0cc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(46),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(11),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(46),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN8_TEMP_1_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10554\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN8_TEMP_0_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10553\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_20_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbf8cbc83b380b08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10062\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(20),
datae => \GRLFPC2_0.FPO.FRAC\(36),
datad => \GRLFPC2_0.FPO.FRAC\(37),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bf838cb0bc808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10064\,
dataf => \GRLFPC2_0.FPO.FRAC\(38),
datae => \GRLFPC2_0.FPO.FRAC\(39),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333ff3ff000cc0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(34),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(23),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(35),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9988\,
dataf => \GRLFPC2_0.FPI.LDOP_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(150),
datac => N_715);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10108\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9988\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_35_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33f33fff00c00ccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(35),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(22),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(35),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_35_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9987\,
dataf => \GRLFPC2_0.FPI.LDOP_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(151),
datac => N_714);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_35_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10107\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(35),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9987\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9991\,
dataf => \GRLFPC2_0.FPI.LDOP_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(147),
datac => N_718);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10111\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(31),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9991\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3fcf0ff030c000")
port map (
combout => N_59331,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(31),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f000f0ffff0ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(31),
dataf => N_59331,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9974\,
dataf => \GRLFPC2_0.FPI.LDOP_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(164),
datac => N_701);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10094\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(48),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9974\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3ff333cc0cc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(48),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(9),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcb3b0bf8c83808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10054\,
dataf => \GRLFPC2_0.FPO.FRAC\(29),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(28),
datad => \GRLFPC2_0.FPO.FRAC\(28),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_45_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10037\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(45),
datae => \GRLFPC2_0.FPO.FRAC\(12),
datad => \GRLFPC2_0.FPO.FRAC\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bf838cb0bc808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10078\,
dataf => \GRLFPC2_0.FPO.FRAC\(52),
datae => \GRLFPC2_0.FPO.FRAC\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10135\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10015\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff0ffff0ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(50),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33f33fff00c00ccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(50),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_20_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10002\,
dataf => \GRLFPC2_0.FPI.LDOP_5\,
datae => \GRLFPC2_0.FPI.OP2\(37),
datad => \GRLFPC2_0.FPI.OP2\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(136));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_20_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10122\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(20),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10002\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_20_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33f33fff00c00ccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(20),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(37),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(20),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_21_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10001\,
dataf => \GRLFPC2_0.FPI.LDOP_5\,
datae => \GRLFPC2_0.FPI.OP2\(36),
datad => \GRLFPC2_0.FPI.OP2\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(137));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_21_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10121\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(21),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10001\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfc00f00fff03f30")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9828\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(39),
datae => N_59328,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_20_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcf3f0ff0c03000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(20),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(20),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_21_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33f33fff00c00ccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(21),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(36),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(21),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(22),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3fcf00f030c00")
port map (
combout => N_59328,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(19),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(20),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_42_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9980\,
dataf => \GRLFPC2_0.FPI.LDOP_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(158),
datac => N_707);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_42_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10100\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(42),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9980\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_42_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33f33fff00c00ccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(42),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(15),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(43),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10051\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(31),
datae => \GRLFPC2_0.FPO.FRAC\(26),
datad => \GRLFPC2_0.FPO.FRAC\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_30_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10052\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(30),
datae => \GRLFPC2_0.FPO.FRAC\(27),
datad => \GRLFPC2_0.FPO.FRAC\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10053\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(29),
datae => \GRLFPC2_0.FPO.FRAC\(28),
datad => \GRLFPC2_0.FPO.FRAC\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_40_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9982\,
dataf => \GRLFPC2_0.FPI.LDOP_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(156),
datac => N_709);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_40_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10102\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(40),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9982\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_40_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333ff3ff000cc0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(40),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(41),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(40),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcff3c33c0c3000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(31),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(30),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9990\,
dataf => \GRLFPC2_0.FPI.LDOP_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(148),
datac => N_717);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10110\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9990\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33c30cfc30c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(32),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(30),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f000f0ffff0ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(32),
dataf => N_59318,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10031\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(51),
datae => \GRLFPC2_0.FPO.FRAC\(6),
datad => \GRLFPC2_0.FPO.FRAC\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10035\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(47),
datae => \GRLFPC2_0.FPO.FRAC\(10),
datad => \GRLFPC2_0.FPO.FRAC\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f00cfc03f30fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9791\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10205\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9969\,
dataf => \GRLFPC2_0.FPI.LDOP_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(169),
datac => N_696);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10089\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(53),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9969\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3ff030cf0fc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10207\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(54),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3cf330cf0cc300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(51),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00ffff0f0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(53),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10207\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbf8cbc83b380b08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10063\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(19),
datae => \GRLFPC2_0.FPO.FRAC\(37),
datad => \GRLFPC2_0.FPO.FRAC\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_38_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9984\,
dataf => \GRLFPC2_0.FPI.LDOP_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(154),
datac => N_711);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_38_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10104\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(38),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9984\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_38_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333ff3ff000cc0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(38),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(19),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(39),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcf3f00f0c0300")
port map (
combout => N_59323,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0f000ffffff0ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(0),
dataf => N_59323,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8_I\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10019\,
dataf => \GRLFPC2_0.FPI.LDOP_4\,
datae => \GRLFPC2_0.FPI.OP2\(54),
datad => \GRLFPC2_0.FPI.OP2\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(119));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10139\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10019\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00fff0ff0fffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(54),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333ff3ff000cc0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(54),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9986\,
dataf => \GRLFPC2_0.FPI.LDOP_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(152),
datac => N_713);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10106\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(36),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9986\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcf3c0cf3c33000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(36),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(36),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(35),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f000f0ffff0ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(36),
dataf => N_59319,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffccfcc33300300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(5),
datae => N_59200,
datad => N_59192,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3fcf00f030c00")
port map (
combout => N_59281,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_46_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cc0fffffcc0f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(46),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(46),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datac => N_59251,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_35_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(35),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(37),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datac => N_59253,
datab => N_59275);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccfffff0cc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(8),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datac => N_59270,
datab => N_59269);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccfffff0cc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(36),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(36),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datac => N_59232,
datab => N_59244);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3fcf0ff030c000")
port map (
combout => N_59319,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(36),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(37),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3fcf00f030c00")
port map (
combout => N_59318,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(33),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_30_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9992\,
dataf => \GRLFPC2_0.FPI.LDOP_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(146),
datac => N_719);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_30_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10112\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(30),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9992\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_30_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcf3f00f0c0300")
port map (
combout => N_59317,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(31),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_30_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffccfcc33300300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(30),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(28),
datae => N_59185,
datad => N_59205,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_30_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3cf330cf0cc300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(30),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(28),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(30),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_30_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f00fff00f0fffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(30),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(30),
datae => N_59317,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10030\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(52),
datae => \GRLFPC2_0.FPO.FRAC\(5),
datad => \GRLFPC2_0.FPO.FRAC\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10136\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10016\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccfffff0cc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datac => N_59265,
datab => N_59264);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8_I\(57),
datad => N_59194,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00fff0ff0fffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(51),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333ff3ff000cc0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(51),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_CIN_2_RNIHRRR7_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c33c3cc33cc3c33c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_60.Z_1_CO1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1281_I\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_58\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.CIN_2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bcb0bf838c808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10079\,
dataf => \GRLFPC2_0.FPO.FRAC\(54),
datae => \GRLFPC2_0.FPO.FRAC\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10018\,
dataf => \GRLFPC2_0.FPI.LDOP_4\,
datae => \GRLFPC2_0.FPI.OP2\(53),
datad => \GRLFPC2_0.FPI.OP2\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(120));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10138\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10018\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccfffff0cc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datac => N_59269,
datab => N_59267);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff0ffff0ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33f33fff00c00ccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(53),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10017\,
dataf => \GRLFPC2_0.FPI.LDOP_4\,
datae => \GRLFPC2_0.FPI.OP2\(52),
datad => \GRLFPC2_0.FPI.OP2\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(121));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10137\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10017\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datac => N_59269,
datab => N_59267);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datac => N_59264,
datab => N_59228);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(5),
dataf => N_59164,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8_I\(57),
datad => N_59200,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00fff0ff0fffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(52),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33f33fff00c00ccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(52),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3fcf00f030c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8_I\(57),
datae => N_59200,
datad => N_59164,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3fcf00f030c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8_I\(57),
datae => N_59194,
datad => N_59163,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_39_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10043\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(39),
datae => \GRLFPC2_0.FPO.FRAC\(18),
datad => \GRLFPC2_0.FPO.FRAC\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_38_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10044\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(38),
datae => \GRLFPC2_0.FPO.FRAC\(19),
datad => \GRLFPC2_0.FPO.FRAC\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10034\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(48),
datae => \GRLFPC2_0.FPO.FRAC\(9),
datad => \GRLFPC2_0.FPO.FRAC\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10028\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(54),
datae => \GRLFPC2_0.FPO.FRAC\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30cf3fc000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6583\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_258_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00fff00ff00fff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8_0\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1281_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_58\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7035\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_4_0_RNIR1HC1_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f3cc3f000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7034\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6961\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bf838cb0bc808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10081\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_176__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_175__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"d9c85140fbea7362")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10027\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_252_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfffcf00c0ffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10530\,
dataf => \GRLFPC2_0.FPO.EXP\(6),
datae => \GRLFPC2_0.FPO.EXP\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(239));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33fc30cf03cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(34),
dataf => N_59205,
datae => N_59172,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_45_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcf3f00f0c0300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(45),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(44),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(43),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10029\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(53),
datae => \GRLFPC2_0.FPO.FRAC\(4),
datad => \GRLFPC2_0.FPO.FRAC\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bcb0bf838c808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10069\,
dataf => \GRLFPC2_0.FPO.FRAC\(44),
datae => \GRLFPC2_0.FPO.FRAC\(43),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_12_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bf838cb0bc808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10070\,
dataf => \GRLFPC2_0.FPO.FRAC\(44),
datae => \GRLFPC2_0.FPO.FRAC\(45),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bf838cb0bc808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10057\,
dataf => \GRLFPC2_0.FPO.FRAC\(31),
datae => \GRLFPC2_0.FPO.FRAC\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN2_DIVMULTV_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000f0000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_DIVMULTV\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_24_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bf838cb0bc808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10058\,
dataf => \GRLFPC2_0.FPO.FRAC\(32),
datae => \GRLFPC2_0.FPO.FRAC\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(24),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10011\,
dataf => \GRLFPC2_0.FPI.LDOP_5\,
datae => \GRLFPC2_0.FPI.OP2\(46),
datad => \GRLFPC2_0.FPI.OP2\(43),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(127));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10131\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(11),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10011\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33f33fff00c00ccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(11),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(46),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bcb0bf838c808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10065\,
dataf => \GRLFPC2_0.FPO.FRAC\(40),
datae => \GRLFPC2_0.FPO.FRAC\(39),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_16_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bf838cb0bc808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10066\,
dataf => \GRLFPC2_0.FPO.FRAC\(40),
datae => \GRLFPC2_0.FPO.FRAC\(41),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_14_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10008\,
dataf => \GRLFPC2_0.FPI.LDOP_5\,
datae => \GRLFPC2_0.FPI.OP2\(43),
datad => \GRLFPC2_0.FPI.OP2\(40),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(130));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_14_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10128\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(14),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10008\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_14_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33f33fff00c00ccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(14),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(43),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(14),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_41_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10041\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(41),
datae => \GRLFPC2_0.FPO.FRAC\(16),
datad => \GRLFPC2_0.FPO.FRAC\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_37_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10045\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(37),
datae => \GRLFPC2_0.FPO.FRAC\(20),
datad => \GRLFPC2_0.FPO.FRAC\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10046\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(36),
datae => \GRLFPC2_0.FPO.FRAC\(21),
datad => \GRLFPC2_0.FPO.FRAC\(20),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_35_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10047\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(35),
datae => \GRLFPC2_0.FPO.FRAC\(22),
datad => \GRLFPC2_0.FPO.FRAC\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10049\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(33),
datae => \GRLFPC2_0.FPO.FRAC\(24),
datad => \GRLFPC2_0.FPO.FRAC\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10050\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(32),
datae => \GRLFPC2_0.FPO.FRAC\(25),
datad => \GRLFPC2_0.FPO.FRAC\(24),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_40_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10042\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(40),
datae => \GRLFPC2_0.FPO.FRAC\(17),
datad => \GRLFPC2_0.FPO.FRAC\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_37_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9985\,
dataf => \GRLFPC2_0.FPI.LDOP_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(153),
datac => N_712);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_37_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10105\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(37),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9985\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_38_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(38),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(40),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datac => N_59232,
datab => N_59244);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_37_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3fcf00f030c00")
port map (
combout => N_59311,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(38),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(37),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_35_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffccfcc33300300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(35),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(33),
datae => N_59218,
datad => N_59197,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(36),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(36),
datae => N_59205,
datad => N_59172,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_37_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3cfc33c300c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(37),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(36),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(35),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(37),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_37_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f00fff00f0fffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(37),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(37),
datae => N_59311,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_41_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9981\,
dataf => \GRLFPC2_0.FPI.LDOP_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(157),
datac => N_708);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_41_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10101\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(41),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9981\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_42_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccfffff0cc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(42),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(42),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datac => N_59251,
datab => N_59249);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_41_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ffffccf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(41),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(41),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datac => N_59254,
datab => N_59255);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_41_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33f33fff00c00ccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(41),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(16),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(41),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN38_SHDVAR_4: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN38_SHDVAR_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03ff03ff000003ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_2_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN17_SHDVAR\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_4\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_2_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333f00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_2_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_2_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_0_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(57),
dataf => N_59189,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3fcf00f030c00")
port map (
combout => N_59229,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(56),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bf838cb0bc808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10071\,
dataf => \GRLFPC2_0.FPO.FRAC\(45),
datae => \GRLFPC2_0.FPO.FRAC\(46),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_0_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_21_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbf8cbc83b380b08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10061\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(21),
datae => \GRLFPC2_0.FPO.FRAC\(35),
datad => \GRLFPC2_0.FPO.FRAC\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_23_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcc00ccf0f0f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9999\,
dataf => \GRLFPC2_0.FPI.LDOP_5\,
datae => \GRLFPC2_0.FPI.OP2\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(139),
datab => N_726);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_23_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10119\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(23),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9999\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_23_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333ff3ff000cc0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(23),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(24),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_22_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10000\,
dataf => \GRLFPC2_0.FPI.LDOP_5\,
datae => \GRLFPC2_0.FPI.OP2\(35),
datad => \GRLFPC2_0.FPI.OP2\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(138));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_22_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10120\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(22),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10000\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_23_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccfffff0cc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(23),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(23),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datac => N_59235,
datab => N_59234);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_22_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccfffff0cc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(22),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(22),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datac => N_59239,
datab => N_59260);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_22_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333ff3ff000cc0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(22),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(35),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(23),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(22),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_22_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3fcf0ff030c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(22),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(22),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(21),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfc0fff00f003f30")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9844\,
dataf => N_59304,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccfffff0cc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datac => N_59264,
datab => N_59228);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59268,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ccf0ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datae => N_59268,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59267,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcf3f00f0c0300")
port map (
combout => N_59304,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffff0000f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8_I\(57),
datae => N_59164,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffff0000f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8_I\(57),
datae => N_59163,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff0ffff0ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(55),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_24_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcc00ccf0f0f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9998\,
dataf => \GRLFPC2_0.FPI.LDOP_5\,
datae => \GRLFPC2_0.FPI.OP2\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(140),
datab => N_725);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_24_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10118\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(24),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9998\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_24_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(24),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(26),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datac => N_59239,
datab => N_59260);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_22_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(22),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(22),
datae => N_59219,
datad => N_59170,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_23_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3fcf00f030c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(23),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(22),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(23),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_24_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333ff3ff000cc0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(24),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(33),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(24),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_22_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bf838cb0bc808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10060\,
dataf => \GRLFPC2_0.FPO.FRAC\(34),
datae => \GRLFPC2_0.FPO.FRAC\(35),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(22),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9995\,
dataf => \GRLFPC2_0.FPI.LDOP_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(143),
datac => N_722);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10115\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(27),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9995\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333ff3ff000cc0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(27),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(30),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(28),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_43_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9979\,
dataf => \GRLFPC2_0.FPI.LDOP_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(159),
datac => N_706);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_43_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10099\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(43),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9979\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_43_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffccf00000ccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(43),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(45),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datac => N_59254,
datab => N_59255);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_41_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcffccc33033000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(41),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(39),
datae => N_59168,
datad => N_59169,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_43_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333ff3ff000cc0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(43),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(14),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(43),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9996\,
dataf => \GRLFPC2_0.FPI.LDOP_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(142),
datac => N_723);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10116\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(26),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9996\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ffffccf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(27),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(27),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datac => N_59235,
datab => N_59236);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333ff3ff000cc0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(26),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(31),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff30f03fcf00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10206\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(54),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffccfcc33300300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(51),
datae => N_59188,
datad => N_59189,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3cfc33c300c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(54),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(53),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00ffff0f0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(54),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(54),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10206\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9968\,
dataf => \GRLFPC2_0.FPI.LDOP_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(170),
datac => N_695);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10088\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(54),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9968\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcc00ccf0f0f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9997\,
dataf => \GRLFPC2_0.FPI.LDOP_5\,
datae => \GRLFPC2_0.FPI.OP2\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(141),
datab => N_724);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10117\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(25),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9997\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9970\,
dataf => \GRLFPC2_0.FPI.LDOP_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(168),
datac => N_697);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10090\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(52),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9970\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9971\,
dataf => \GRLFPC2_0.FPI.LDOP_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(167),
datac => N_698);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10091\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(51),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9971\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9972\,
dataf => \GRLFPC2_0.FPI.LDOP_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(166),
datac => N_699);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10092\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(50),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9972\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_39_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9983\,
dataf => \GRLFPC2_0.FPI.LDOP_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(155),
datac => N_710);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_39_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10103\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(39),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9983\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9994\,
dataf => \GRLFPC2_0.FPI.LDOP_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(144),
datac => N_721);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10114\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(28),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9994\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0ffc0cf303f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10208\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(54),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(53),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3fcc0cf333c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(52),
dataf => N_59211,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(52),
datad => N_59210,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3cfc33c300c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(52),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(51),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(50),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00ffff0f0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(52),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(52),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10208\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcf3f0ff0c03000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10209\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(51),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(51),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(51),
datae => N_59186,
datad => N_59188,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3ccf0cf330c300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(51),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(51),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(49),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ffff0f000f0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(51),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10209\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ffffccf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(51),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(51),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcf3f00f0c0300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10210\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(51),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcffccc33033000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(50),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(48),
datae => N_59211,
datad => N_59210,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(50),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(49),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(49),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00ffff0f0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(50),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(50),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10210\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_15_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59232,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_14_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59254,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_39_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3fcf0ff030c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(39),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(39),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(38),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_22_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59197,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_37_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(37),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(37),
datae => N_59218,
datad => N_59197,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_23_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59172,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_38_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3fcf00f030c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(38),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(37),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(38),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_39_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33f33fff00c00ccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(39),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(18),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(39),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(40),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffccf00000ccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(28),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(30),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datac => N_59239,
datab => N_59240);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(26),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(26),
datae => N_59170,
datad => N_59171,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33f33fff00c00ccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(28),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(29),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(28),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffccf00000ccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(29),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(31),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datac => N_59235,
datab => N_59236);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcf3f0ff0c03000")
port map (
combout => N_59309,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(29),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3fcc0cf333c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(29),
dataf => N_59213,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(29),
datad => N_59166,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcffccc33033000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(27),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(25),
datae => N_59213,
datad => N_59166,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3cfc33c300c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(29),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(28),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f000f0ffff0ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(29),
dataf => N_59309,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9993\,
dataf => \GRLFPC2_0.FPI.LDOP_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(145),
datac => N_720);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10113\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(29),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9993\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffcc0f0000cc0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(48),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(50),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datac => N_59251,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cc0fffffcc0f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(47),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(47),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datac => N_59252,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_46_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcf3f0ff0c03000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(46),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(46),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(43),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(47),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(10),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9975\,
dataf => \GRLFPC2_0.FPI.LDOP_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(163),
datac => N_702);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10095\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(47),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9975\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_14_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffccf00000ccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(14),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(16),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datac => N_59270,
datab => N_59271);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => N_59308,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(14),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0cc00ccffcc0fcc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9833\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(44),
datae => N_59308,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfc00f00fff03f30")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9790\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(1),
datae => N_59297,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(114),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10003\,
dataf => \GRLFPC2_0.FPI.LDOP_5\,
datae => \GRLFPC2_0.FPI.OP2\(38),
datad => \GRLFPC2_0.FPI.OP2\(35),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(135));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10123\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(19),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10003\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59196,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(56),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(56),
datae => N_59211,
datad => N_59195,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59211,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59195,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffc3330cfcc0300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(54),
dataf => N_59211,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(52),
datad => N_59195,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59189,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(55),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(55),
datae => N_59188,
datad => N_59189,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(19),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(21),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datac => N_59272,
datab => N_59263);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcf3f00f0c0300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(19),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(18),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3fcc0cf333c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(18),
dataf => N_59219,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(18),
datad => N_59183,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3fcf0ff030c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(18),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(18),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333ff3ff000cc0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(19),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(38),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(20),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_20_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33fc30cf03cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(20),
dataf => N_59219,
datae => N_59170,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_21_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3fcf00f030c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(21),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(20),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(21),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59240,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59239,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59245,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ffffccf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(26),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(26),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datac => N_59239,
datab => N_59240);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59274,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_30_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59273,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59235,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59234,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(25),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(27),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datac => N_59235,
datab => N_59234);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59179,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_21_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccfffff0cc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(21),
dataf => N_59179,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_35_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59220,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_22_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccfffff0cc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(22),
dataf => N_59220,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_37_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59170,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59171,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_24_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffccfcc33300300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(24),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(22),
datae => N_59170,
datad => N_59171,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_24_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3fcf0ff030c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(24),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(24),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(23),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333ff3ff000cc0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(25),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(26),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_81_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0ff00ccccff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(81),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => N_694,
datac => N_665,
datab => N_601);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_80_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ffccfff000cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(80),
dataf => \GRLFPC2_0.FPI.OP1\(32),
datae => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_666,
datab => N_602);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_10_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bcb0bf838c808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10072\,
dataf => \GRLFPC2_0.FPO.FRAC\(47),
datae => \GRLFPC2_0.FPO.FRAC\(46),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_77_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ffcc00f000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(77),
dataf => \GRLFPC2_0.FPI.OP1\(38),
datae => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_666,
datab => N_602);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_74_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ffccfff000cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(74),
dataf => \GRLFPC2_0.FPI.OP1\(38),
datae => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_672,
datab => N_608);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_71_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ffcc00f000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(71),
dataf => \GRLFPC2_0.FPI.OP1\(44),
datae => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_672,
datab => N_608);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_65_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ffccfff000cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(65),
dataf => \GRLFPC2_0.FPI.OP1\(47),
datae => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_681,
datab => N_617);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ffcc00f000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(62),
dataf => \GRLFPC2_0.FPI.OP1\(53),
datae => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_681,
datab => N_617);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_78_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ffcc00f000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(78),
dataf => \GRLFPC2_0.FPI.OP1\(37),
datae => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_665,
datab => N_601);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_75_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ffccfff000cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(75),
dataf => \GRLFPC2_0.FPI.OP1\(37),
datae => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_671,
datab => N_607);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_72_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ffcc00f000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(72),
dataf => \GRLFPC2_0.FPI.OP1\(43),
datae => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_671,
datab => N_607);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_69_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ffccfff000cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(69),
dataf => \GRLFPC2_0.FPI.OP1\(43),
datae => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_677,
datab => N_613);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_66_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ffcc00f000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(66),
dataf => \GRLFPC2_0.FPI.OP1\(49),
datae => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_677,
datab => N_613);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_41_254_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ffccfff000cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_41\(254),
dataf => \GRLFPC2_0.FPI.OP1\(55),
datae => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_689,
datab => N_625);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_76_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ffccfff000cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(76),
dataf => \GRLFPC2_0.FPI.OP1\(36),
datae => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_670,
datab => N_606);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_73_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ffcc00f000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(73),
dataf => \GRLFPC2_0.FPI.OP1\(42),
datae => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_670,
datab => N_606);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_70_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ffccfff000cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(70),
dataf => \GRLFPC2_0.FPI.OP1\(42),
datae => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_676,
datab => N_612);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_67_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ffcc00f000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(67),
dataf => \GRLFPC2_0.FPI.OP1\(48),
datae => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_676,
datab => N_612);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ffccfff000cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(61),
dataf => \GRLFPC2_0.FPI.OP1\(51),
datae => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_685,
datab => N_621);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10015\,
dataf => \GRLFPC2_0.FPI.LDOP_5\,
datae => \GRLFPC2_0.FPI.OP2\(50),
datad => \GRLFPC2_0.FPI.OP2\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(123));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bf838cb0bc808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10077\,
dataf => \GRLFPC2_0.FPO.FRAC\(51),
datae => \GRLFPC2_0.FPO.FRAC\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_12_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10010\,
dataf => \GRLFPC2_0.FPI.LDOP_5\,
datae => \GRLFPC2_0.FPI.OP2\(45),
datad => \GRLFPC2_0.FPI.OP2\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(128));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_12_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10130\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(12),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10010\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccfffff0cc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(13),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(13),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datac => N_59263,
datab => N_59262);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_12_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ffffccf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(12),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(12),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datac => N_59270,
datab => N_59271);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_12_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3ccc03f330c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(12),
dataf => N_59191,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(12),
datad => N_59217,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_12_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3fcf0ff030c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(12),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(12),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_10_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffccfcc33300300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(10),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(8),
datae => N_59191,
datad => N_59217,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_12_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33f33fff00c00ccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(12),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(45),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(12),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_16_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0ff000cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10006\,
dataf => \GRLFPC2_0.FPI.LDOP_5\,
datae => \GRLFPC2_0.FPI.OP2\(38),
datad => \GRLFPC2_0.FPI.OP2\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(132));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_16_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10126\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(16),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10006\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_15_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10007\,
dataf => \GRLFPC2_0.FPI.LDOP_5\,
datae => \GRLFPC2_0.FPI.OP2\(42),
datad => \GRLFPC2_0.FPI.OP2\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(131));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_15_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10127\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(15),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10007\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_16_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffc0f0cf3f00300")
port map (
combout => N_59294,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(18),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_16_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcff3c33c0c3000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(16),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(15),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(16),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(14),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_16_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f00fff00f0fffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(16),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(16),
datae => N_59294,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_15_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcff0c03f0f3000")
port map (
combout => N_59293,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(18),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(15),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_15_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3ccf0cf330c300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(15),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(15),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(14),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_15_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f00fff00f0fffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(15),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(15),
datae => N_59293,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10048\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(34),
datae => \GRLFPC2_0.FPO.FRAC\(23),
datad => \GRLFPC2_0.FPO.FRAC\(22),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_49_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ccf0cc0fccffcc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9797\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10211\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_49_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffcc0f0000cc0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(49),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(51),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datac => N_59252,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_49_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcf3f0ff0c03000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10211\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(49),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59188,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_49_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffccfcc33300300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(49),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(47),
datae => N_59186,
datad => N_59188,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_49_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcf3f0ff0c03000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(49),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(49),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(46),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_12_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59186,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_10_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59187,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59210,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcf3f00f0c0300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(48),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(47),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(46),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_44_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9978\,
dataf => \GRLFPC2_0.FPI.LDOP_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(160),
datac => N_705);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_44_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10098\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(44),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9978\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_10_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59255,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59252,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_12_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59250,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_9_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59251,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59249,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_44_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0ccfffff0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(44),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(46),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datac => N_59251,
datab => N_59249);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_44_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3ff333cc0cc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(44),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(44),
datae => N_59209,
datad => N_59208,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_21_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59206,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59208,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_15_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59209,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_42_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcffccc33033000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(42),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(40),
datae => N_59209,
datad => N_59208,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_20_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59169,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_16_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59168,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59199,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_43_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3ff333cc0cc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(43),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(43),
datae => N_59168,
datad => N_59169,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_44_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33f33fff00c00ccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(44),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(13),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10032\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(50),
datae => \GRLFPC2_0.FPO.FRAC\(7),
datad => \GRLFPC2_0.FPO.FRAC\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_49_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10033\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(49),
datae => \GRLFPC2_0.FPO.FRAC\(8),
datad => \GRLFPC2_0.FPO.FRAC\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0cc00ccffcc0fcc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9829\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(40),
datae => N_59291,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59260,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_35_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59261,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_39_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59271,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59272,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_38_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59263,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_40_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59246,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3ff030cf0fc000")
port map (
combout => N_59291,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(18),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(20),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(17),
dataf => N_59178,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3fcf00f030c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(17),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(16),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_44_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59178,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_46_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59173,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_15_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(15),
dataf => N_59173,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccff00f0f0f0f0")
port map (
combout => N_59217,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_45_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59183,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_41_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59219,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_16_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcf3303fccc3000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(16),
dataf => N_59219,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(14),
datad => N_59183,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10016\,
dataf => \GRLFPC2_0.FPI.LDOP_4\,
datae => \GRLFPC2_0.FPI.OP2\(51),
datad => \GRLFPC2_0.FPI.OP2\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(122));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9989\,
dataf => \GRLFPC2_0.FPI.LDOP_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(149),
datac => N_716);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10109\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(33),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9989\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59238,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_21_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59243,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59244,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_23_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59242,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59253,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_22_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59275,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_20_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59237,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_24_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59236,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccfffff0cc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(33),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(33),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datac => N_59253,
datab => N_59275);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_24_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59180,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(33),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(33),
datae => N_59213,
datad => N_59218,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59174,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_30_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59213,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59218,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33fc30cf03cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(31),
dataf => N_59213,
datae => N_59218,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59185,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59205,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffccf3c03f0c3300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(32),
dataf => N_59185,
datae => N_59205,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333ff3ff000cc0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(33),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(24),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_116_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_118_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_0_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_122_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21));
\GRLFPC2_0_COMB_DBGDATA_4_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(1),
dataf => \GRLFPC2_0.R.FSR.CEXC\(1),
datae => N_397,
datad => N_398,
datac => N_664,
datab => N_600);
\GRLFPC2_0_COMB_DBGDATA_4_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(3),
dataf => \GRLFPC2_0.R.FSR.CEXC\(3),
datae => N_397,
datad => N_398,
datac => N_666,
datab => N_602);
\GRLFPC2_0_FPI_OP1_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP1\(33),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => N_600,
datad => N_664);
\GRLFPC2_0_FPI_OP1_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP1\(36),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => N_603,
datad => N_667);
\GRLFPC2_0_COMB_WRDATA_4_9_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(9),
dataf => \GRLFPC2_0.R.I.RES\(38),
datae => \GRLFPC2_0.R.I.RES\(9),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_WRDATA_9_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(9),
dataf => N_412,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_372,
datab => \GRLFPC2_0.COMB.WRDATA_4\(9));
\GRLFPC2_0_COMB_WRDATA_4_41_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(41),
dataf => \GRLFPC2_0.R.I.RES\(38),
datae => \GRLFPC2_0.R.I.RES\(41),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_WRDATA_41_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(9),
dataf => N_412,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_372,
datab => \GRLFPC2_0.COMB.WRDATA_4\(41));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_14_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00f0f0ff00cccc")
port map (
combout => \GRLFPC2_0.N_3152\,
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.FSR.FTT\(0),
datac => N_677,
datab => N_613);
\GRLFPC2_0_FPI_OP2_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(55),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_654,
datad => N_718);
\GRLFPC2_0_FPI_OP2_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(56),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_655,
datad => N_719);
\GRLFPC2_0_FPI_OP2_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(58),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_657,
datad => N_721);
\GRLFPC2_0_FPI_OP2_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(59),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_658,
datad => N_722);
\GRLFPC2_0_FPI_OP2_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(60),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_659,
datad => N_723);
\GRLFPC2_0_FPI_OP2_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(61),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_660,
datad => N_724);
\GRLFPC2_0_FPI_OP2_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(62),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_661,
datad => N_725);
\GRLFPC2_0_COMB_DBGDATA_4_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(25),
dataf => \GRLFPC2_0.R.FSR.TEM\(2),
datae => N_397,
datad => N_398,
datac => N_688,
datab => N_624);
\GRLFPC2_0_RS1_1_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => RFI2_RD1ADDRZ(0),
dataf => \GRLFPC2_0.COMB.RS1_1\(1),
datae => N_399,
datad => N_395);
\GRLFPC2_0_RS1_1_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => RFI2_RD1ADDRZ(1),
dataf => \GRLFPC2_0.COMB.RS1_1\(2),
datae => N_400,
datad => N_395);
\GRLFPC2_0_RS1_1_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => RFI2_RD1ADDRZ(2),
dataf => \GRLFPC2_0.COMB.RS1_1\(3),
datae => N_401,
datad => N_395);
\GRLFPC2_0_RS1_1_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => RFI2_RD1ADDRZ(3),
dataf => \GRLFPC2_0.COMB.RS1_1\(4),
datae => N_402,
datad => N_395);
\GRLFPC2_0_RS2_1_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => RFI2_RD2ADDRZ(0),
dataf => \GRLFPC2_0.COMB.RS2_1\(1),
datae => N_399,
datad => N_395);
\GRLFPC2_0_RS2_1_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => RFI2_RD2ADDRZ(1),
dataf => \GRLFPC2_0.COMB.RS2_1\(2),
datae => N_400,
datad => N_395);
\GRLFPC2_0_RS2_1_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => RFI2_RD2ADDRZ(2),
dataf => \GRLFPC2_0.COMB.RS2_1\(3),
datae => N_401,
datad => N_395);
\GRLFPC2_0_RS2_1_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => RFI2_RD2ADDRZ(3),
dataf => \GRLFPC2_0.COMB.RS2_1\(4),
datae => N_402,
datad => N_395);
\GRLFPC2_0_COMB_RF2REN_1_0_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00fcffff00fc0000")
port map (
combout => \GRLFPC2_0.N_3032\,
dataf => \GRLFPC2_0.R.A.RF2REN\(2),
datae => N_9,
datad => \GRLFPC2_0.COMB.LOCKGEN.LOCKI_I_I\,
datac => \GRLFPC2_0.COMB.RS2D_1\,
datab => \GRLFPC2_0.COMB.RS2_1\(0));
\GRLFPC2_0_COMB_RF2REN_1_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0fffffff0ff0000")
port map (
combout => RFI2_REN2Z,
dataf => \GRLFPC2_0.N_3032\,
datae => N_395,
datad => N_396,
datac => N_397);
\GRLFPC2_0_COMB_RF2REN_1_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0fffffff0ff0000")
port map (
combout => RFI2_REN1Z,
dataf => \GRLFPC2_0.N_3033\,
datae => N_395,
datad => N_396,
datac => N_397);
\GRLFPC2_0_COMB_RF1REN_1_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0fffffff0ff0000")
port map (
combout => RFI1_REN2Z,
dataf => \GRLFPC2_0.N_3226\,
datae => N_395,
datad => N_396,
datac => N_397);
\GRLFPC2_0_COMB_RF1REN_1_0_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f300fffff3000000")
port map (
combout => \GRLFPC2_0.N_3227\,
dataf => \GRLFPC2_0.R.A.RF1REN\(1),
datae => N_9,
datad => \GRLFPC2_0.COMB.V.A.RF2REN_1_1\(1),
datac => \GRLFPC2_0.COMB.RS1D_1\,
datab => \GRLFPC2_0.COMB.RS1_1\(0));
\GRLFPC2_0_COMB_RF1REN_1_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0fffffff0ff0000")
port map (
combout => RFI1_REN1Z,
dataf => \GRLFPC2_0.N_3227\,
datae => N_395,
datad => N_396,
datac => N_397);
\GRLFPC2_0_FPI_OP2_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(32),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_631,
datad => N_695);
\GRLFPC2_0_FPI_OP2_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(33),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_632,
datad => N_696);
\GRLFPC2_0_FPI_OP2_49_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(49),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_648,
datad => N_712);
\GRLFPC2_0_FPI_OP2_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(50),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_649,
datad => N_713);
\GRLFPC2_0_FPI_OP2_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(51),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_650,
datad => N_714);
\GRLFPC2_0_FPI_OP2_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(52),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_651,
datad => N_715);
\GRLFPC2_0_FPI_OP2_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(53),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_652,
datad => N_716);
\GRLFPC2_0_FPI_OP2_41_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(41),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_640,
datad => N_704);
\GRLFPC2_0_FPI_OP2_42_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(42),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_641,
datad => N_705);
\GRLFPC2_0_FPI_OP2_43_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(43),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_642,
datad => N_706);
\GRLFPC2_0_FPI_OP2_44_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(44),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_643,
datad => N_707);
\GRLFPC2_0_FPI_OP2_46_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(46),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_645,
datad => N_709);
\GRLFPC2_0_FPI_OP2_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(47),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_646,
datad => N_710);
\GRLFPC2_0_FPI_OP2_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(34),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_633,
datad => N_697);
\GRLFPC2_0_FPI_OP2_35_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(35),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_634,
datad => N_698);
\GRLFPC2_0_FPI_OP2_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(36),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_635,
datad => N_699);
\GRLFPC2_0_FPI_OP2_37_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(37),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_636,
datad => N_700);
\GRLFPC2_0_FPI_OP2_38_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(38),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_637,
datad => N_701);
\GRLFPC2_0_FPI_OP2_39_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(39),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_638,
datad => N_702);
\GRLFPC2_0_FPI_OP2_40_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(40),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_639,
datad => N_703);
\GRLFPC2_0_FPI_OP1_49_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP1\(49),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => N_616,
datad => N_680);
\GRLFPC2_0_COMB_DBGDATA_4_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(13),
dataf => \GRLFPC2_0.N_835\,
datae => N_397,
datad => N_398,
datac => N_676,
datab => N_612);
\GRLFPC2_0_COMB_DBGDATA_4_16_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(16),
dataf => \GRLFPC2_0.R.FSR.FTT\(2),
datae => N_397,
datad => N_398,
datac => N_679,
datab => N_615);
\GRLFPC2_0_FPI_OP1_44_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP1\(44),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => N_611,
datad => N_675);
\GRLFPC2_0_COMB_DBGDATA_4_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(27),
dataf => \GRLFPC2_0.R.FSR.TEM\(4),
datae => N_397,
datad => N_398,
datac => N_690,
datab => N_626);
\GRLFPC2_0_FPI_OP1_38_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP1\(38),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => N_605,
datad => N_669);
\GRLFPC2_0_COMB_V_E_STDATA_1_1_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00f0f0ff00cccc")
port map (
combout => \GRLFPC2_0.N_3146\,
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.FSR.AEXC\(3),
datac => N_671,
datab => N_607);
\GRLFPC2_0_COMB_V_E_STDATA_1_1_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00f0f0ff00cccc")
port map (
combout => \GRLFPC2_0.N_3145\,
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.FSR.AEXC\(2),
datac => N_670,
datab => N_606);
\GRLFPC2_0_COMB_DBGDATA_4_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(6),
dataf => \GRLFPC2_0.R.FSR.AEXC\(1),
datae => N_397,
datad => N_398,
datac => N_669,
datab => N_605);
\GRLFPC2_0_COMB_WRDATA_4_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(36),
dataf => \GRLFPC2_0.R.I.RES\(33),
datae => \GRLFPC2_0.R.I.RES\(36),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_WRDATA_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(4),
dataf => N_407,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_367,
datab => \GRLFPC2_0.COMB.WRDATA_4\(36));
\GRLFPC2_0_WRADDR_1_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRADDRZ(0),
dataf => N_399,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.WRADDR_1_SQMUXA\,
datac => \GRLFPC2_0.R.I.INST\(26),
datab => N_352);
\GRLFPC2_0_WRADDR_1_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRADDRZ(1),
dataf => N_400,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.WRADDR_1_SQMUXA\,
datac => \GRLFPC2_0.R.I.INST\(27),
datab => N_353);
\GRLFPC2_0_WRADDR_1_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRADDRZ(3),
dataf => N_402,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.WRADDR_1_SQMUXA\,
datac => \GRLFPC2_0.R.I.INST\(29),
datab => N_355);
\GRLFPC2_0_COMB_V_I_PC_1_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.R.I.PC\(27),
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.PC_O\(27),
datad => \GRLFPC2_0.FPCI_O\(310));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33cc00f3f3c0c0")
port map (
combout => \GRLFPC2_0.N_3134\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.INST\(29),
datad => \GRLFPC2_0.FPCI_O\(312),
datac => \GRLFPC2_0.R.I.PC_O\(29),
datab => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_COMB_V_E_STDATA_1_0_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33cc00f3f3c0c0")
port map (
combout => \GRLFPC2_0.N_3136\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.INST\(31),
datad => \GRLFPC2_0.FPCI_O\(314),
datac => \GRLFPC2_0.R.I.PC_O\(31),
datab => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_COMB_V_E_STDATA_1_1_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00f0f0ff00cccc")
port map (
combout => \GRLFPC2_0.N_3151\,
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.N_835\,
datac => N_676,
datab => N_612);
\GRLFPC2_0_WRDATA_43_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(11),
dataf => N_414,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_374,
datab => \GRLFPC2_0.COMB.WRDATA_4\(43));
\GRLFPC2_0_FPI_OP1_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP1\(47),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => N_614,
datad => N_678);
\GRLFPC2_0_FPI_OP1_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP1\(52),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => N_619,
datad => N_683);
\GRLFPC2_0_COMB_DBGDATA_4_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(0),
dataf => \GRLFPC2_0.R.FSR.CEXC\(0),
datae => N_397,
datad => N_398,
datac => N_663,
datab => N_599);
\GRLFPC2_0_COMB_DBGDATA_4_9_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(9),
dataf => \GRLFPC2_0.R.FSR.AEXC\(4),
datae => N_397,
datad => N_398,
datac => N_672,
datab => N_608);
\GRLFPC2_0_FPI_OP1_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP1\(32),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => N_599,
datad => N_663);
\GRLFPC2_0_COMB_V_E_STDATA_1_1_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00f0f0ff00cccc")
port map (
combout => \GRLFPC2_0.N_3140\,
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.FSR.CEXC\(2),
datac => N_665,
datab => N_601);
\GRLFPC2_0_FPI_OP1_37_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP1\(37),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => N_604,
datad => N_668);
\GRLFPC2_0_COMB_V_E_STDATA_1_1_9_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00f0f0ff00cccc")
port map (
combout => \GRLFPC2_0.N_3147\,
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.FSR.AEXC\(4),
datac => N_672,
datab => N_608);
\GRLFPC2_0_FPI_OP1_42_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP1\(42),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => N_609,
datad => N_673);
\GRLFPC2_0_FPI_OP1_43_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP1\(43),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => N_610,
datad => N_674);
\GRLFPC2_0_FPI_OP1_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP1\(48),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => N_615,
datad => N_679);
\GRLFPC2_0_COMB_V_E_STDATA_1_1_22_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00f0f0ff00cccc")
port map (
combout => \GRLFPC2_0.N_3160\,
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.FSR.NONSTD\,
datac => N_685,
datab => N_621);
\GRLFPC2_0_WRDATA_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(8),
dataf => N_411,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_371,
datab => \GRLFPC2_0.COMB.WRDATA_4\(8));
\GRLFPC2_0_COMB_WRDATA_4_40_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(40),
dataf => \GRLFPC2_0.R.I.RES\(37),
datae => \GRLFPC2_0.R.I.RES\(40),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_WRDATA_40_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(8),
dataf => N_411,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_371,
datab => \GRLFPC2_0.COMB.WRDATA_4\(40));
\GRLFPC2_0_WRDATA_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(1),
dataf => N_404,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_364,
datab => \GRLFPC2_0.COMB.WRDATA_4\(1));
\GRLFPC2_0_WRDATA_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(5),
dataf => N_408,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_368,
datab => \GRLFPC2_0.COMB.WRDATA_4\(5));
\GRLFPC2_0_COMB_WRDATA_4_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(7),
dataf => \GRLFPC2_0.R.I.RES\(36),
datae => \GRLFPC2_0.R.I.RES\(7),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_WRDATA_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(7),
dataf => N_410,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_370,
datab => \GRLFPC2_0.COMB.WRDATA_4\(7));
\GRLFPC2_0_WRDATA_24_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(24),
dataf => N_427,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_387,
datab => \GRLFPC2_0.COMB.WRDATA_4\(24));
\GRLFPC2_0_WRDATA_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(26),
dataf => N_429,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_389,
datab => \GRLFPC2_0.COMB.WRDATA_4\(26));
\GRLFPC2_0_WRDATA_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(27),
dataf => N_430,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_390,
datab => \GRLFPC2_0.COMB.WRDATA_4\(27));
\GRLFPC2_0_WRDATA_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(29),
dataf => N_432,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_392,
datab => \GRLFPC2_0.COMB.WRDATA_4\(29));
\GRLFPC2_0_COMB_WRDATA_4_30_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(30),
dataf => \GRLFPC2_0.R.I.RES\(59),
datae => \GRLFPC2_0.R.I.RES\(30),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_WRDATA_30_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(30),
dataf => N_433,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_393,
datab => \GRLFPC2_0.COMB.WRDATA_4\(30));
\GRLFPC2_0_COMB_WRDATA_4_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(31),
dataf => \GRLFPC2_0.R.I.RES\(63),
datae => \GRLFPC2_0.R.I.RES\(31),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_WRDATA_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(31),
dataf => N_434,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_394,
datab => \GRLFPC2_0.COMB.WRDATA_4\(31));
\GRLFPC2_0_COMB_WRDATA_4_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(33),
dataf => \GRLFPC2_0.R.I.RES\(30),
datae => \GRLFPC2_0.R.I.RES\(33),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_WRDATA_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(1),
dataf => N_404,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_364,
datab => \GRLFPC2_0.COMB.WRDATA_4\(33));
\GRLFPC2_0_WRDATA_37_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(5),
dataf => N_408,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_368,
datab => \GRLFPC2_0.COMB.WRDATA_4\(37));
\GRLFPC2_0_COMB_WRDATA_4_39_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(39),
dataf => \GRLFPC2_0.R.I.RES\(36),
datae => \GRLFPC2_0.R.I.RES\(39),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_WRDATA_39_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(7),
dataf => N_410,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_370,
datab => \GRLFPC2_0.COMB.WRDATA_4\(39));
\GRLFPC2_0_WRDATA_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(24),
dataf => N_427,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_387,
datab => \GRLFPC2_0.COMB.WRDATA_4\(56));
\GRLFPC2_0_WRDATA_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(26),
dataf => N_429,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_389,
datab => \GRLFPC2_0.COMB.WRDATA_4\(58));
\GRLFPC2_0_WRDATA_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(27),
dataf => N_430,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_390,
datab => \GRLFPC2_0.COMB.WRDATA_4\(59));
\GRLFPC2_0_COMB_WRDATA_4_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(61),
dataf => \GRLFPC2_0.R.I.RES\(58),
datae => \GRLFPC2_0.R.I.RES\(61),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_WRDATA_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(29),
dataf => N_432,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_392,
datab => \GRLFPC2_0.COMB.WRDATA_4\(61));
\GRLFPC2_0_WRDATA_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(30),
dataf => N_433,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_393,
datab => \GRLFPC2_0.COMB.WRDATA_4\(62));
\GRLFPC2_0_WRDATA_63_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(31),
dataf => N_434,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_394,
datab => \GRLFPC2_0.R.I.RES\(63));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33cc00f3f3c0c0")
port map (
combout => \GRLFPC2_0.N_3122\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.INST\(17),
datad => \GRLFPC2_0.FPCI_O\(300),
datac => \GRLFPC2_0.R.I.PC_O\(17),
datab => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_COMB_V_I_PC_1_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.R.I.PC\(18),
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.PC_O\(18),
datad => \GRLFPC2_0.FPCI_O\(301));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_20_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33cc00f3f3c0c0")
port map (
combout => \GRLFPC2_0.N_3125\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.INST\(20),
datad => \GRLFPC2_0.FPCI_O\(303),
datac => \GRLFPC2_0.R.I.PC_O\(20),
datab => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_COMB_V_I_PC_1_24_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.R.I.PC\(24),
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.PC_O\(24),
datad => \GRLFPC2_0.FPCI_O\(307));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_I_M2_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33cc00f3f3c0c0")
port map (
combout => \GRLFPC2_0.N_145\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.INST\(4),
datad => \GRLFPC2_0.FPCI_O\(287),
datac => \GRLFPC2_0.R.I.PC_O\(4),
datab => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_COMB_V_E_STDATA_1_0_I_M2_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33cc00f3f3c0c0")
port map (
combout => \GRLFPC2_0.N_146\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.INST\(5),
datad => \GRLFPC2_0.FPCI_O\(288),
datac => \GRLFPC2_0.R.I.PC_O\(5),
datab => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_COMB_V_I_PC_1_I_M2_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.N_3426\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.PC_O\(6),
datad => \GRLFPC2_0.FPCI_O\(289));
\GRLFPC2_0_COMB_V_I_PC_1_I_M2_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.N_3427\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.PC_O\(7),
datad => \GRLFPC2_0.FPCI_O\(290));
\GRLFPC2_0_COMB_V_I_PC_1_I_M2_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.N_3428\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.PC_O\(8),
datad => \GRLFPC2_0.FPCI_O\(291));
\GRLFPC2_0_COMB_V_I_PC_1_I_M2_9_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.N_3429\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.PC_O\(9),
datad => \GRLFPC2_0.FPCI_O\(292));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_I_M2_10_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33cc00f3f3c0c0")
port map (
combout => \GRLFPC2_0.N_151\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.INST\(10),
datad => \GRLFPC2_0.FPCI_O\(293),
datac => \GRLFPC2_0.R.I.PC_O\(10),
datab => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_COMB_V_E_STDATA_1_0_I_M2_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33cc00f3f3c0c0")
port map (
combout => \GRLFPC2_0.N_152\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.INST\(11),
datad => \GRLFPC2_0.FPCI_O\(294),
datac => \GRLFPC2_0.R.I.PC_O\(11),
datab => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_COMB_V_E_STDATA_1_0_I_M2_12_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33cc00f3f3c0c0")
port map (
combout => \GRLFPC2_0.N_153\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.INST\(12),
datad => \GRLFPC2_0.FPCI_O\(295),
datac => \GRLFPC2_0.R.I.PC_O\(12),
datab => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_COMB_V_I_PC_1_I_M2_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.N_140\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.PC_O\(13),
datad => \GRLFPC2_0.FPCI_O\(296));
\GRLFPC2_0_COMB_V_I_PC_1_I_M2_14_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.N_141\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.PC_O\(14),
datad => \GRLFPC2_0.FPCI_O\(297));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_I_M2_15_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33cc00f3f3c0c0")
port map (
combout => \GRLFPC2_0.N_156\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.INST\(15),
datad => \GRLFPC2_0.FPCI_O\(298),
datac => \GRLFPC2_0.R.I.PC_O\(15),
datab => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_COMB_V_E_STDATA_1_0_I_M2_16_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33cc00f3f3c0c0")
port map (
combout => \GRLFPC2_0.N_157\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.INST\(16),
datad => \GRLFPC2_0.FPCI_O\(299),
datac => \GRLFPC2_0.R.I.PC_O\(16),
datab => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_COMB_DBGDATA_4_23_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(23),
dataf => \GRLFPC2_0.R.FSR.TEM\(0),
datae => N_397,
datad => N_398,
datac => N_686,
datab => N_622);
\GRLFPC2_0_COMB_DBGDATA_4_24_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(24),
dataf => \GRLFPC2_0.R.FSR.TEM\(1),
datae => N_397,
datad => N_398,
datac => N_687,
datab => N_623);
\GRLFPC2_0_COMB_DBGDATA_4_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(31),
dataf => \GRLFPC2_0.R.FSR.RD\(1),
datae => N_397,
datad => N_398,
datac => N_694,
datab => N_630);
\GRLFPC2_0_FPI_OP1_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP1\(55),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => N_622,
datad => N_686);
\GRLFPC2_0_COMB_WRDATA_4_22_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(22),
dataf => \GRLFPC2_0.R.I.RES\(51),
datae => \GRLFPC2_0.R.I.RES\(22),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_WRDATA_22_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(22),
dataf => N_425,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_385,
datab => \GRLFPC2_0.COMB.WRDATA_4\(22));
\GRLFPC2_0_WRDATA_23_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(23),
dataf => N_426,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_386,
datab => \GRLFPC2_0.COMB.WRDATA_4\(23));
\GRLFPC2_0_COMB_WRDATA_4_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(54),
dataf => \GRLFPC2_0.R.I.RES\(51),
datae => \GRLFPC2_0.R.I.RES\(54),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_WRDATA_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(22),
dataf => N_425,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_385,
datab => \GRLFPC2_0.COMB.WRDATA_4\(54));
\GRLFPC2_0_WRDATA_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(23),
dataf => N_426,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_386,
datab => \GRLFPC2_0.COMB.WRDATA_4\(55));
\GRLFPC2_0_COMB_WRDATA_4_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(26),
dataf => \GRLFPC2_0.R.I.RES\(55),
datae => \GRLFPC2_0.R.I.RES\(26),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_DBGDATA_4_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(26),
dataf => \GRLFPC2_0.R.FSR.TEM\(3),
datae => N_397,
datad => N_398,
datac => N_689,
datab => N_625);
\GRLFPC2_0_COMB_V_E_STDATA_1_1_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00f0f0ff00cccc")
port map (
combout => \GRLFPC2_0.N_3164\,
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.FSR.TEM\(3),
datac => N_689,
datab => N_625);
\GRLFPC2_0_WRDATA_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(0),
dataf => N_403,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_363,
datab => \GRLFPC2_0.COMB.WRDATA_4\(0));
\GRLFPC2_0_WRDATA_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(2),
dataf => N_405,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_365,
datab => \GRLFPC2_0.COMB.WRDATA_4\(2));
\GRLFPC2_0_WRDATA_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(11),
dataf => N_414,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_374,
datab => \GRLFPC2_0.COMB.WRDATA_4\(11));
\GRLFPC2_0_COMB_WRDATA_4_14_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(14),
dataf => \GRLFPC2_0.R.I.RES\(43),
datae => \GRLFPC2_0.R.I.RES\(14),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_WRDATA_14_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(14),
dataf => N_417,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_377,
datab => \GRLFPC2_0.COMB.WRDATA_4\(14));
\GRLFPC2_0_WRDATA_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(17),
dataf => N_420,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_380,
datab => \GRLFPC2_0.COMB.WRDATA_4\(17));
\GRLFPC2_0_COMB_WRDATA_4_20_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(20),
dataf => \GRLFPC2_0.R.I.RES\(49),
datae => \GRLFPC2_0.R.I.RES\(20),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_WRDATA_20_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(20),
dataf => N_423,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_383,
datab => \GRLFPC2_0.COMB.WRDATA_4\(20));
\GRLFPC2_0_WRDATA_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(0),
dataf => N_403,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_363,
datab => \GRLFPC2_0.COMB.WRDATA_4\(32));
\GRLFPC2_0_WRDATA_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(2),
dataf => N_405,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_365,
datab => \GRLFPC2_0.COMB.WRDATA_4\(34));
\GRLFPC2_0_WRDATA_46_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(14),
dataf => N_417,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_377,
datab => \GRLFPC2_0.COMB.WRDATA_4\(46));
\GRLFPC2_0_WRDATA_49_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(17),
dataf => N_420,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_380,
datab => \GRLFPC2_0.COMB.WRDATA_4\(49));
\GRLFPC2_0_WRDATA_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(20),
dataf => N_423,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_383,
datab => \GRLFPC2_0.COMB.WRDATA_4\(52));
\GRLFPC2_0_COMB_DBGDATA_4_22_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(22),
dataf => \GRLFPC2_0.R.FSR.NONSTD\,
datae => N_397,
datad => N_398,
datac => N_685,
datab => N_621);
\GRLFPC2_0_WRDATA_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(13),
dataf => N_416,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_376,
datab => \GRLFPC2_0.COMB.WRDATA_4\(13));
\GRLFPC2_0_WRDATA_16_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(16),
dataf => N_419,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_379,
datab => \GRLFPC2_0.COMB.WRDATA_4\(16));
\GRLFPC2_0_WRDATA_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(19),
dataf => N_422,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_382,
datab => \GRLFPC2_0.COMB.WRDATA_4\(19));
\GRLFPC2_0_WRDATA_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(25),
dataf => N_428,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_388,
datab => \GRLFPC2_0.COMB.WRDATA_4\(25));
\GRLFPC2_0_WRDATA_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(28),
dataf => N_431,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_391,
datab => \GRLFPC2_0.COMB.WRDATA_4\(28));
\GRLFPC2_0_WRDATA_45_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(13),
dataf => N_416,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_376,
datab => \GRLFPC2_0.COMB.WRDATA_4\(45));
\GRLFPC2_0_WRDATA_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(16),
dataf => N_419,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_379,
datab => \GRLFPC2_0.COMB.WRDATA_4\(48));
\GRLFPC2_0_WRDATA_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(19),
dataf => N_422,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_382,
datab => \GRLFPC2_0.COMB.WRDATA_4\(51));
\GRLFPC2_0_WRDATA_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(25),
dataf => N_428,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_388,
datab => \GRLFPC2_0.COMB.WRDATA_4\(57));
\GRLFPC2_0_COMB_WRDATA_4_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(60),
dataf => \GRLFPC2_0.R.I.RES\(57),
datae => \GRLFPC2_0.R.I.RES\(60),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_WRDATA_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(28),
dataf => N_431,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_391,
datab => \GRLFPC2_0.COMB.WRDATA_4\(60));
\GRLFPC2_0_WRDATA_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(3),
dataf => N_406,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_366,
datab => \GRLFPC2_0.COMB.WRDATA_4\(3));
\GRLFPC2_0_COMB_WRDATA_4_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(6),
dataf => \GRLFPC2_0.R.I.RES\(35),
datae => \GRLFPC2_0.R.I.RES\(6),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_WRDATA_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(6),
dataf => N_409,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_369,
datab => \GRLFPC2_0.COMB.WRDATA_4\(6));
\GRLFPC2_0_COMB_WRDATA_4_12_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(12),
dataf => \GRLFPC2_0.R.I.RES\(41),
datae => \GRLFPC2_0.R.I.RES\(12),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_WRDATA_12_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(12),
dataf => N_415,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_375,
datab => \GRLFPC2_0.COMB.WRDATA_4\(12));
\GRLFPC2_0_COMB_WRDATA_4_15_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(15),
dataf => \GRLFPC2_0.R.I.RES\(44),
datae => \GRLFPC2_0.R.I.RES\(15),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_WRDATA_15_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(15),
dataf => N_418,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_378,
datab => \GRLFPC2_0.COMB.WRDATA_4\(15));
\GRLFPC2_0_COMB_WRDATA_4_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(18),
dataf => \GRLFPC2_0.R.I.RES\(47),
datae => \GRLFPC2_0.R.I.RES\(18),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_WRDATA_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(18),
dataf => N_421,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_381,
datab => \GRLFPC2_0.COMB.WRDATA_4\(18));
\GRLFPC2_0_COMB_WRDATA_4_21_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(21),
dataf => \GRLFPC2_0.R.I.RES\(50),
datae => \GRLFPC2_0.R.I.RES\(21),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_WRDATA_21_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(21),
dataf => N_424,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_384,
datab => \GRLFPC2_0.COMB.WRDATA_4\(21));
\GRLFPC2_0_WRDATA_35_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(3),
dataf => N_406,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_366,
datab => \GRLFPC2_0.COMB.WRDATA_4\(35));
\GRLFPC2_0_COMB_WRDATA_4_38_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(38),
dataf => \GRLFPC2_0.R.I.RES\(35),
datae => \GRLFPC2_0.R.I.RES\(38),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_WRDATA_38_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(6),
dataf => N_409,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_369,
datab => \GRLFPC2_0.COMB.WRDATA_4\(38));
\GRLFPC2_0_COMB_WRDATA_4_44_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(44),
dataf => \GRLFPC2_0.R.I.RES\(41),
datae => \GRLFPC2_0.R.I.RES\(44),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_WRDATA_44_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(12),
dataf => N_415,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_375,
datab => \GRLFPC2_0.COMB.WRDATA_4\(44));
\GRLFPC2_0_COMB_WRDATA_4_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(47),
dataf => \GRLFPC2_0.R.I.RES\(44),
datae => \GRLFPC2_0.R.I.RES\(47),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_WRDATA_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(15),
dataf => N_418,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_378,
datab => \GRLFPC2_0.COMB.WRDATA_4\(47));
\GRLFPC2_0_COMB_WRDATA_4_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(50),
dataf => \GRLFPC2_0.R.I.RES\(47),
datae => \GRLFPC2_0.R.I.RES\(50),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_WRDATA_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(18),
dataf => N_421,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_381,
datab => \GRLFPC2_0.COMB.WRDATA_4\(50));
\GRLFPC2_0_COMB_WRDATA_4_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(53),
dataf => \GRLFPC2_0.R.I.RES\(50),
datae => \GRLFPC2_0.R.I.RES\(53),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_WRDATA_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(21),
dataf => N_424,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_384,
datab => \GRLFPC2_0.COMB.WRDATA_4\(53));
\GRLFPC2_0_COMB_V_I_PC_1_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.R.I.PC\(2),
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.PC_O\(2),
datad => \GRLFPC2_0.FPCI_O\(285));
\GRLFPC2_0_COMB_V_I_PC_1_21_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.R.I.PC\(21),
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.PC_O\(21),
datad => \GRLFPC2_0.FPCI_O\(304));
\GRLFPC2_0_COMB_V_I_PC_1_22_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.R.I.PC\(22),
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.PC_O\(22),
datad => \GRLFPC2_0.FPCI_O\(305));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_23_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33cc00f3f3c0c0")
port map (
combout => \GRLFPC2_0.N_3128\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.INST\(23),
datad => \GRLFPC2_0.FPCI_O\(306),
datac => \GRLFPC2_0.R.I.PC_O\(23),
datab => \GRLFPC2_0.COMB.V.E.STDATA2\);
\GRLFPC2_0_COMB_V_I_PC_1_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.R.I.PC\(26),
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.PC_O\(26),
datad => \GRLFPC2_0.FPCI_O\(309));
\GRLFPC2_0_WRDATA_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(4),
dataf => N_407,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_367,
datab => \GRLFPC2_0.COMB.WRDATA_4\(4));
\GRLFPC2_0_WRDATA_42_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(10),
dataf => N_413,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_373,
datab => \GRLFPC2_0.COMB.WRDATA_4\(42));
\GRLFPC2_0_COMB_WRDATA_4_43_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(43),
dataf => \GRLFPC2_0.R.I.RES\(40),
datae => \GRLFPC2_0.R.I.RES\(43),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(8),
dataf => \GRLFPC2_0.R.I.RES\(37),
datae => \GRLFPC2_0.R.I.RES\(8),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(1),
dataf => \GRLFPC2_0.R.I.RES\(30),
datae => \GRLFPC2_0.R.I.RES\(1),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(5),
dataf => \GRLFPC2_0.R.I.RES\(34),
datae => \GRLFPC2_0.R.I.RES\(5),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_24_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(24),
dataf => \GRLFPC2_0.R.I.RES\(53),
datae => \GRLFPC2_0.R.I.RES\(24),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(27),
dataf => \GRLFPC2_0.R.I.RES\(56),
datae => \GRLFPC2_0.R.I.RES\(27),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(29),
dataf => \GRLFPC2_0.R.I.RES\(58),
datae => \GRLFPC2_0.R.I.RES\(29),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_37_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(37),
dataf => \GRLFPC2_0.R.I.RES\(34),
datae => \GRLFPC2_0.R.I.RES\(37),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(56),
dataf => \GRLFPC2_0.R.I.RES\(53),
datae => \GRLFPC2_0.R.I.RES\(56),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(58),
dataf => \GRLFPC2_0.R.I.RES\(55),
datae => \GRLFPC2_0.R.I.RES\(58),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(59),
dataf => \GRLFPC2_0.R.I.RES\(56),
datae => \GRLFPC2_0.R.I.RES\(59),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(62),
dataf => \GRLFPC2_0.R.I.RES\(59),
datae => \GRLFPC2_0.R.I.RES\(62),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_23_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(23),
dataf => \GRLFPC2_0.R.I.RES\(52),
datae => \GRLFPC2_0.R.I.RES\(23),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(55),
dataf => \GRLFPC2_0.R.I.RES\(52),
datae => \GRLFPC2_0.R.I.RES\(55),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(0),
dataf => \GRLFPC2_0.R.I.RES\(29),
datae => \GRLFPC2_0.R.I.RES\(0),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(2),
dataf => \GRLFPC2_0.R.I.RES\(31),
datae => \GRLFPC2_0.R.I.RES\(2),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(11),
dataf => \GRLFPC2_0.R.I.RES\(40),
datae => \GRLFPC2_0.R.I.RES\(11),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(17),
dataf => \GRLFPC2_0.R.I.RES\(46),
datae => \GRLFPC2_0.R.I.RES\(17),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(32),
dataf => \GRLFPC2_0.R.I.RES\(29),
datae => \GRLFPC2_0.R.I.RES\(32),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(34),
dataf => \GRLFPC2_0.R.I.RES\(31),
datae => \GRLFPC2_0.R.I.RES\(34),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_46_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(46),
dataf => \GRLFPC2_0.R.I.RES\(43),
datae => \GRLFPC2_0.R.I.RES\(46),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_49_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(49),
dataf => \GRLFPC2_0.R.I.RES\(46),
datae => \GRLFPC2_0.R.I.RES\(49),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(52),
dataf => \GRLFPC2_0.R.I.RES\(49),
datae => \GRLFPC2_0.R.I.RES\(52),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(13),
dataf => \GRLFPC2_0.R.I.RES\(42),
datae => \GRLFPC2_0.R.I.RES\(13),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_16_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(16),
dataf => \GRLFPC2_0.R.I.RES\(45),
datae => \GRLFPC2_0.R.I.RES\(16),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(19),
dataf => \GRLFPC2_0.R.I.RES\(48),
datae => \GRLFPC2_0.R.I.RES\(19),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(25),
dataf => \GRLFPC2_0.R.I.RES\(54),
datae => \GRLFPC2_0.R.I.RES\(25),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(28),
dataf => \GRLFPC2_0.R.I.RES\(57),
datae => \GRLFPC2_0.R.I.RES\(28),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_45_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(45),
dataf => \GRLFPC2_0.R.I.RES\(42),
datae => \GRLFPC2_0.R.I.RES\(45),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(48),
dataf => \GRLFPC2_0.R.I.RES\(45),
datae => \GRLFPC2_0.R.I.RES\(48),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(51),
dataf => \GRLFPC2_0.R.I.RES\(48),
datae => \GRLFPC2_0.R.I.RES\(51),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(57),
dataf => \GRLFPC2_0.R.I.RES\(54),
datae => \GRLFPC2_0.R.I.RES\(57),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(3),
dataf => \GRLFPC2_0.R.I.RES\(32),
datae => \GRLFPC2_0.R.I.RES\(3),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_35_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(35),
dataf => \GRLFPC2_0.R.I.RES\(32),
datae => \GRLFPC2_0.R.I.RES\(35),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(4),
dataf => \GRLFPC2_0.R.I.RES\(33),
datae => \GRLFPC2_0.R.I.RES\(4),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_COMB_WRDATA_4_42_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(42),
dataf => \GRLFPC2_0.R.I.RES\(39),
datae => \GRLFPC2_0.R.I.RES\(42),
datad => \GRLFPC2_0.COMB.RDD_2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_2_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00fc30ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_2_RNI51QB6_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cf0000fc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(375),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_15: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_15\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_22: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000300000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_22\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_15\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_26: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000003f00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_26\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_22\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_20: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_20\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_19: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_19\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_17: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_17\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_23: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000300000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_23\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_17\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_27: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0003000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_27\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_23\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_19\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_112_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(112),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(112),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(112));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_111_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(111),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(111),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(111));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_110_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(110),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(110),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(110));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_109_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(109),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(109),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(109));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_108_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(108),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(108),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(108));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_107_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(107),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(107),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(107));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_102_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(102),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(102),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(102));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_96_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(96),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(96),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(96));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_93_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(93),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(93),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(93));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_79_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(79),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_70_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(70),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(70),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(70));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_67_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(67),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(67),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(67));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_66_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(66),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(66),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(66));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_64_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(64),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(64),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(64));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(62),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(62),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(62));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_113_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaff00f0f0cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(113),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_106_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaff00f0f0cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(106),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datad => \GRLFPC2_0.FPO.FRAC\(9),
datac => \GRLFPC2_0.FPO.FRAC\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_105_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaff00f0f0cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(105),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datad => \GRLFPC2_0.FPO.FRAC\(10),
datac => \GRLFPC2_0.FPO.FRAC\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_104_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaff00f0f0cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(104),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datad => \GRLFPC2_0.FPO.FRAC\(11),
datac => \GRLFPC2_0.FPO.FRAC\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_103_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaff00f0f0cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(103),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datad => \GRLFPC2_0.FPO.FRAC\(12),
datac => \GRLFPC2_0.FPO.FRAC\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_86_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaff00f0f0cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(86),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datad => \GRLFPC2_0.FPO.FRAC\(29),
datac => \GRLFPC2_0.FPO.FRAC\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_85_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaff00f0f0cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(85),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datad => \GRLFPC2_0.FPO.FRAC\(30),
datac => \GRLFPC2_0.FPO.FRAC\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_84_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaff00f0f0cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(84),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datad => \GRLFPC2_0.FPO.FRAC\(31),
datac => \GRLFPC2_0.FPO.FRAC\(29),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_81_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaff00f0f0cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(81),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(34),
datac => \GRLFPC2_0.FPO.FRAC\(32),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_80_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaff00f0f0cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(80),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(35),
datac => \GRLFPC2_0.FPO.FRAC\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_79_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccff00f0f0aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(79),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(36),
datac => \GRLFPC2_0.FPO.FRAC\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_70_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccff00f0f0aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(70),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(45),
datac => \GRLFPC2_0.FPO.FRAC\(43),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_67_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccff00f0f0aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(67),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(48),
datac => \GRLFPC2_0.FPO.FRAC\(46),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_66_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccff00f0f0aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(66),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(49),
datac => \GRLFPC2_0.FPO.FRAC\(47),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_64_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccff00f0f0aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(64),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(51),
datac => \GRLFPC2_0.FPO.FRAC\(49),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccf0f0ff00aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(62),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(51),
datac => \GRLFPC2_0.FPO.FRAC\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaff00f0f0cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(58),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_176__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_115_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(115),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(115));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_114_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(114),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(114));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNISVH7OR2_29_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(29),
dataf => N_26534,
datae => N_26536,
datad => N_26535);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIH8IFPR2_30_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(30),
dataf => N_26534,
datae => N_26538,
datad => N_26537);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_RNIOQOJ0S2_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(31),
dataf => N_26534,
datae => N_26540,
datad => N_26539);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNISMK1AS2_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(32),
dataf => N_26534,
datae => N_26542,
datad => N_26541);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI8FCTSS2_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(33),
dataf => N_26534,
datae => N_26544,
datad => N_26543);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI40SK2U2_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(34),
dataf => N_26534,
datae => N_26546,
datad => N_26545);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI02R3E03_35_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(35),
dataf => N_26534,
datae => N_26548,
datad => N_26547);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIS5P1553_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(36),
dataf => N_26534,
datae => N_26550,
datad => N_26549);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIODLTIE3_37_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(37),
dataf => N_26534,
datae => N_26552,
datad => N_26551);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIKTDLE1_38_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(38),
dataf => N_26534,
datae => N_26554,
datad => N_26553);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIGTU4671_39_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(39),
dataf => N_26534,
datae => N_26556,
datad => N_26555);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIGC14LI3_40_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(40),
dataf => N_26534,
datae => N_26558,
datad => N_26557);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIKA62J9_41_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(41),
dataf => N_26534,
datae => N_26560,
datad => N_26559);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIKLQALP1_45_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(45),
dataf => N_26534,
datae => N_26568,
datad => N_26567);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIGTOFJN_46_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(46),
dataf => N_26534,
datae => N_26570,
datad => N_26569);
\GRLFPC2_0_WRDATA_10_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(10),
dataf => N_413,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_373,
datab => \GRLFPC2_0.COMB.WRDATA_4\(10));
GRLFPC2_0_COMB_WREN2_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffc000000fc00")
port map (
combout => RFI2_WRENZ,
dataf => N_398,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => N_9,
datac => \GRLFPC2_0.COMB.WREN2_9_IV_1\,
datab => \GRLFPC2_0.COMB.WREN2_9_IV_0\);
\GRLFPC2_0_WRADDR_1_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRADDRZ(2),
dataf => N_401,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.WRADDR_1_SQMUXA\,
datac => \GRLFPC2_0.R.I.INST\(28),
datab => N_354);
GRLFPC2_0_COMB_WREN1_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000fc00fffffc00")
port map (
combout => RFI1_WRENZ,
dataf => N_398,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => N_9,
datac => \GRLFPC2_0.COMB.WREN1_9_IV_1\,
datab => \GRLFPC2_0.COMB.WREN1_9_IV_0\);
\GRLFPC2_0_COMB_V_I_PC_1_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.R.I.PC\(28),
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.PC_O\(28),
datad => \GRLFPC2_0.FPCI_O\(311));
\GRLFPC2_0_COMB_V_I_PC_1_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.R.I.PC\(25),
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.PC_O\(25),
datad => \GRLFPC2_0.FPCI_O\(308));
\GRLFPC2_0_COMB_WRDATA_4_10_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(10),
dataf => \GRLFPC2_0.R.I.RES\(39),
datae => \GRLFPC2_0.R.I.RES\(10),
datad => \GRLFPC2_0.COMB.RDD_2\);
GRLFPC2_0_COMB_WREN2_9_IV_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffc00fc00fc00")
port map (
combout => \GRLFPC2_0.COMB.WREN2_9_IV_1\,
dataf => \GRLFPC2_0.WREN2_2_SQMUXA\,
datae => N_351,
datad => \GRLFPC2_0.WREN2_1_SQMUXA_0\,
datac => N_359,
datab => N_358);
GRLFPC2_0_COMB_WREN2_9_IV_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000f0cc0000")
port map (
combout => \GRLFPC2_0.COMB.WREN2_9_IV_0\,
dataf => \GRLFPC2_0.COMB.RDD_2\,
datae => \GRLFPC2_0.N_1586\,
datad => \GRLFPC2_0.WRADDR_1_SQMUXA\,
datac => \GRLFPC2_0.R.I.INST\(25),
datab => N_351);
GRLFPC2_0_WREN1_1_SQMUXA_1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000003000000000")
port map (
combout => \GRLFPC2_0.WREN2_1_SQMUXA_0\,
dataf => N_346,
datae => \GRLFPC2_0.R.X.SEQERR\,
datad => \GRLFPC2_0.N_1105\,
datac => \GRLFPC2_0.R.X.LD\,
datab => \GRLFPC2_0.R.X.AFSR\);
GRLFPC2_0_COMB_WREN1_9_IV_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300ffff03000300")
port map (
combout => \GRLFPC2_0.COMB.WREN1_9_IV_1\,
dataf => \GRLFPC2_0.WREN2_2_SQMUXA\,
datae => N_351,
datad => \GRLFPC2_0.WREN2_1_SQMUXA_0\,
datac => N_359,
datab => N_358);
GRLFPC2_0_COMB_WREN1_9_IV_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00000f330000")
port map (
combout => \GRLFPC2_0.COMB.WREN1_9_IV_0\,
dataf => \GRLFPC2_0.COMB.RDD_2\,
datae => \GRLFPC2_0.N_1586\,
datad => \GRLFPC2_0.WRADDR_1_SQMUXA\,
datac => \GRLFPC2_0.R.I.INST\(25),
datab => N_351);
\GRLFPC2_0_FPI_OP1_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP1\(60),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => N_627,
datad => N_691);
GRLFPC2_0_WREN2_2_SQMUXA: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000030")
port map (
combout => \GRLFPC2_0.WREN2_2_SQMUXA\,
dataf => \GRLFPC2_0.N_1105\,
datae => N_346,
datad => \GRLFPC2_0.R.X.SEQERR\,
datac => \GRLFPC2_0.R.X.LD\,
datab => \GRLFPC2_0.R.X.AFSR\);
GRLFPC2_0_R_I_V_ENA_RNO_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff0f")
port map (
combout => \GRLFPC2_0.R.I.V_1_0_G0_I_O4_2\,
dataf => \GRLFPC2_0.N_1570\,
datae => \GRLFPC2_0.N_1470\,
datad => \GRLFPC2_0.COMB.ANNULRES_1\,
datac => N_7);
GRLFPC2_0_COMB_UN3_HOLDN: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0000")
port map (
combout => \GRLFPC2_0.N_1237\,
dataf => N_154,
datae => N_153);
GRLFPC2_0_COMB_UN1_FPCI_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0000")
port map (
combout => \GRLFPC2_0.N_1683\,
dataf => N_223,
datae => N_222);
GRLFPC2_0_ANNULRES_0_SQMUXA_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000c0")
port map (
combout => \GRLFPC2_0.N_1676\,
dataf => \GRLFPC2_0.R.X.FPOP\,
datae => \GRLFPC2_0.R.I.EXEC\,
datad => \GRLFPC2_0.R.M.FPOP\,
datac => \GRLFPC2_0.R.E.FPOP\,
datab => \GRLFPC2_0.N_1683\);
GRLFPC2_0_ANNULFPU_0_SQMUXA_0_A3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000000000")
port map (
combout => \GRLFPC2_0.N_1675_1\,
dataf => \GRLFPC2_0.R.M.FPOP\,
datae => N_291,
datad => N_292);
GRLFPC2_0_R_I_V_ENA_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f000f000f00030")
port map (
combout => \GRLFPC2_0.R.I.V_1_0_G2\,
dataf => \GRLFPC2_0.N_1255\,
datae => \GRLFPC2_0.N_1470\,
datad => \GRLFPC2_0.COMB.ANNULRES_1\,
datac => N_7,
datab => N_9);
GRLFPC2_0_R_I_V_ENA: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffc000cffff0000")
port map (
combout => N_48775,
dataf => \GRLFPC2_0.V.FSR.CEXC_3_SQMUXA_1\,
datae => \GRLFPC2_0.R.I.V_1_0_G2\,
datad => \GRLFPC2_0.N_1255\,
datac => \GRLFPC2_0.R.I.V_1_0_G0_I_O4_2\,
datab => \GRLFPC2_0.R.I.V\);
\GRLFPC2_0_COMB_V_I_PC_1_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.R.I.PC\(3),
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.PC_O\(3),
datad => \GRLFPC2_0.FPCI_O\(286));
\GRLFPC2_0_COMB_DBGDATA_4_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(2),
dataf => \GRLFPC2_0.R.FSR.CEXC\(2),
datae => N_397,
datad => N_398,
datac => N_665,
datab => N_601);
\GRLFPC2_0_COMB_V_E_STDATA_1_1_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00f0f0ff00cccc")
port map (
combout => \GRLFPC2_0.N_3141\,
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.FSR.CEXC\(3),
datac => N_666,
datab => N_602);
\GRLFPC2_0_COMB_DBGDATA_4_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(4),
dataf => \GRLFPC2_0.R.FSR.CEXC\(4),
datae => N_397,
datad => N_398,
datac => N_667,
datab => N_603);
\GRLFPC2_0_R_FSR_FCC_RNO_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfc0cfc0cfcfc0c0")
port map (
combout => \GRLFPC2_0.R.FSR.FCC_0_0_0__G1\,
dataf => \GRLFPC2_0.N_1515\,
datae => \GRLFPC2_0.N_3219\,
datad => \GRLFPC2_0.R.I.CC\(0),
datac => \GRLFPC2_0.N_1517\,
datab => N_413);
\GRLFPC2_0_R_FSR_FCC_RNO_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfc0cfc0cfcfc0c0")
port map (
combout => \GRLFPC2_0.R.FSR.FCC_0_0_1__G1\,
dataf => \GRLFPC2_0.N_1515\,
datae => \GRLFPC2_0.N_3220\,
datad => \GRLFPC2_0.R.I.CC\(1),
datac => \GRLFPC2_0.N_1517\,
datab => N_414);
\GRLFPC2_0_COMB_V_A_RF1REN_1_1_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.COMB.V.A.RF2REN_1_1\(1),
dataf => \GRLFPC2_0.COMB.LOCKGEN.LOCKI_I_I\,
datae => \GRLFPC2_0.COMB.RS1V_1\);
\GRLFPC2_0_FPI_OP1_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP1\(57),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => N_624,
datad => N_688);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_41_255_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ffcc00f000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_41\(255),
dataf => \GRLFPC2_0.FPI.OP1\(57),
datae => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_685,
datab => N_621);
\GRLFPC2_0_FPI_OP1_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP1\(61),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => N_628,
datad => N_692);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_41_251_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ffcc00f000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_41\(251),
dataf => \GRLFPC2_0.FPI.OP1\(61),
datae => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_689,
datab => N_625);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_251_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10517\,
dataf => \GRLFPC2_0.FPO.EXP\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(238));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_255_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10513\,
dataf => \GRLFPC2_0.FPO.EXP\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242));
\GRLFPC2_0_FPI_OP1_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP1\(56),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => N_623,
datad => N_687);
\GRLFPC2_0_FPI_OP1_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP1\(53),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => N_620,
datad => N_684);
\GRLFPC2_0_FPI_OP1_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP1\(59),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => N_626,
datad => N_690);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_246_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfffcf00c0ffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10536\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\(12),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_247_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfffcf00c0ffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10535\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\(11),
datae => \GRLFPC2_0.FPO.EXP\(10),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_250_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfffcf00c0ffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10532\,
dataf => \GRLFPC2_0.FPO.EXP\(8),
datae => \GRLFPC2_0.FPO.EXP\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(237));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_256_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfffc0ffcf00c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10526\,
dataf => \GRLFPC2_0.FPO.EXP\(1),
datae => \GRLFPC2_0.FPO.EXP\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(243));
\GRLFPC2_0_FPI_OP2_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(57),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_656,
datad => N_720);
\GRLFPC2_0_FPI_OP2_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(54),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_653,
datad => N_717);
\GRLFPC2_0_COMB_V_STATE_7_IV_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000003cf00cf")
port map (
combout => \GRLFPC2_0.N_1309\,
dataf => \GRLFPC2_0.N_1570\,
datae => \GRLFPC2_0.N_1213\,
datad => \GRLFPC2_0.R.STATE\(0),
datac => \GRLFPC2_0.R.X.SEQERR\,
datab => \GRLFPC2_0.N_1105\);
\GRLFPC2_0_COMB_V_STATE_1_IV_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f000f000c000000")
port map (
combout => \GRLFPC2_0.R.STATE_0_0_1__I0_I_1\,
dataf => \GRLFPC2_0.N_1721\,
datae => CPO_EXCZ,
datad => N_7,
datac => \GRLFPC2_0.N_1669\,
datab => N_11);
\GRLFPC2_0_COMB_DBGDATA_4_30_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(30),
dataf => \GRLFPC2_0.R.FSR.RD\(0),
datae => N_397,
datad => N_398,
datac => N_693,
datab => N_629);
\GRLFPC2_0_FPI_OP1_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP1\(62),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => N_629,
datad => N_693);
\GRLFPC2_0_COMB_V_I_PC_1_30_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.R.I.PC\(30),
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.PC_O\(30),
datad => \GRLFPC2_0.FPCI_O\(313));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN53_SCTRL_NEW: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00030003ff030003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.U_RDN_1\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.UN17_U_RDN\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.TEMP\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_U_RDN_1_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff3f0f3f0f3f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.U_RDN_1\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(21),
datad => \GRLFPC2_0.R.FSR.RD\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SIGNRESULT: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cccc0003c3cc0c")
port map (
combout => \GRLFPC2_0.FPO.SIGN\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(12),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(24),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(23));
\GRLFPC2_0_FPI_OP2_63_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(63),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_662,
datad => N_726);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_2_IV_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"e4f5ffff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_I_I_0\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_IV_0\(0),
datae => N_29788,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4233\,
datac => \GRLFPC2_0.FPO.SIGN\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(22));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_UN17_U_RDN: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f000f000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.UN17_U_RDN\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(21),
datad => \GRLFPC2_0.R.FSR.RD\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59166,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datac => N_59228,
datab => N_59226);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59228,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00f0f0f0f0")
port map (
combout => N_59226,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc30fc30fc30cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10936\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10939\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff00f0f0f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10937\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ccccff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10936\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(243));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff000000ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff000000ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff000000ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIQ83D_43_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10939\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_NORMDETECT_NOTSLFROMNORM_19_0_A2_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00fc00cf00ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M13\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM12\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M12_RNI0U1C_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0f0f00000f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M13\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM12\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M8_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff00ff00ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M8\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M13_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000fff30000fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M13\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M8\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M2_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff0000ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M2\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M12_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000fff30000fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M2\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TEMP\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_64_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff00ff")
port map (
combout => \GRLFPC2_0.FPI.RST\,
dataf => \GRLFPC2_0.R.MK.RST\,
datae => \GRLFPC2_0.R.MK.RST2\,
datad => N_7);
GRLFPC2_0_R_MK_HOLDN1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffffffff")
port map (
combout => \GRLFPC2_0.N_2101\,
dataf => \GRLFPC2_0.R.MK.RST2\,
datae => N_7);
GRLFPC2_0_FPCO_HOLDN_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => CPO_HOLDNZ,
dataf => \GRLFPC2_0.R.MK.HOLDN1\,
datae => \GRLFPC2_0.R.MK.HOLDN2\);
\GRLFPC2_0_COMB_V_E_STDATA_1_0_I_M2_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33cc00f3f3c0c0")
port map (
combout => \GRLFPC2_0.N_158\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.INST\(19),
datad => \GRLFPC2_0.FPCI_O\(302),
datac => \GRLFPC2_0.R.I.PC_O\(19),
datab => \GRLFPC2_0.COMB.V.E.STDATA2\);
GRLFPC2_0_COMB_RDD_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff3fffc0000000")
port map (
combout => \GRLFPC2_0.COMB.RDD_2\,
dataf => \GRLFPC2_0.R.I.RDD\,
datae => \GRLFPC2_0.R.X.RDD\,
datad => \GRLFPC2_0.V.I.EXEC_0_SQMUXA\,
datac => \GRLFPC2_0.R.I.V\,
datab => \GRLFPC2_0.COMB.UN1_R.I.V_1\);
GRLFPC2_0_COMB_QNE2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => \GRLFPC2_0.N_835\,
dataf => \GRLFPC2_0.R.STATE\(1),
datae => \GRLFPC2_0.R.STATE\(0));
\GRLFPC2_0_FPI_OP1_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP1\(51),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => N_618,
datad => N_682);
GRLFPC2_0_ANNULRES_0_SQMUXA_4_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => \GRLFPC2_0.COMB.UN1_R.I.V_1\,
dataf => \GRLFPC2_0.R.X.FPOP\,
datae => \GRLFPC2_0.R.I.EXEC\);
GRLFPC2_0_COMB_UN1_FPCI: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff00")
port map (
combout => \GRLFPC2_0.N_1105\,
dataf => N_10,
datae => N_360,
datad => N_361);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_14_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bf838cb0bc808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10068\,
dataf => \GRLFPC2_0.FPO.FRAC\(42),
datae => \GRLFPC2_0.FPO.FRAC\(43),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(14),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNISV3N6J_43_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(43),
dataf => N_26534,
datae => N_26564,
datad => N_26563);
\GRLFPC2_0_R_I_CC_RNO_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f000f0000000f0")
port map (
combout => \GRLFPC2_0.R.I.CC_0_0_1__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(40),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(39));
\GRLFPC2_0_R_I_CC_RNO_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f000f000f00000")
port map (
combout => \GRLFPC2_0.R.I.CC_0_0_0__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(40),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(39));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_TEMP: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4233\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIG3MJ_40_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4662\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(39),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(38),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(40));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_65_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccff00f0f0aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(65),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(50),
datac => \GRLFPC2_0.FPO.FRAC\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_65_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(65),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(65),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(65));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI07GUEN1_42_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(42),
dataf => N_26534,
datae => N_26562,
datad => N_26561);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_9_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10133\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(9),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10013\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67));
\GRLFPC2_0_FPI_OP2_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(48),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_647,
datad => N_711);
\GRLFPC2_0_FPI_OP2_45_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP2\(45),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => N_644,
datad => N_708);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_9_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10013\,
dataf => \GRLFPC2_0.FPI.LDOP_5\,
datae => \GRLFPC2_0.FPI.OP2\(48),
datad => \GRLFPC2_0.FPI.OP2\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(125));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_41_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59258,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_43_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59270,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59269,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_10_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(10),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(12),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datac => N_59270,
datab => N_59269);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_42_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59262,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_44_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_59265,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_59264,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_9_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(9),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(11),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datac => N_59265,
datab => N_59264);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M8_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M8\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M13_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0f03ffff0f00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M13\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M8\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIOHB8MA2_44_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(44),
dataf => N_26534,
datae => N_26566,
datad => N_26565);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\(8),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccff00f0f0f0f0")
port map (
combout => N_59191,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(240));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccff00f0f0f0f0")
port map (
combout => N_59194,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(238));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_49_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccff00f0f0f0f0")
port map (
combout => N_59193,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccf0f0ff00ff00")
port map (
combout => N_59200,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(237));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccff00f0f0f0f0")
port map (
combout => N_59192,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(241));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(239));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ccf0ffff0000")
port map (
combout => N_59215,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(243));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_9_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(9),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(9),
datae => N_59200,
datad => N_59192,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_9_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3fcf0ff030c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(9),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(9),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M12_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f0000000c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M2\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M14S2_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M2_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M2\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN25_GEN: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c0c000c000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN25_GEN\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SCLSBS_2\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SCLSBS_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_954\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7210\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN2_MIXOIN_3_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff00f0f0f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_3_I\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.NOTPROP_3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN25_GEN\,
datac => N_59288);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN2_MIXOIN_2_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcffc0fc00c000")
port map (
combout => N_59288,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SBLSBS_1\(1),
datae => N_59286,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_959_I\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SBLSBS_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5452\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_0_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_NOTPROP: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0cfcfffff3f3ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.NOTPROP\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10579\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5322\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(371));
GRLFPC2_0_COMB_RS2D_1_IV: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0c0c000c0c0000")
port map (
combout => \GRLFPC2_0.COMB.RS2D_1\,
dataf => \GRLFPC2_0.COMB.FPDECODE.RS1D5\,
datae => \GRLFPC2_0.N_896\,
datad => \GRLFPC2_0.N_884\,
datac => N_80,
datab => N_81);
GRLFPC2_0_RS1D_CNST_0_O2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0c00000000f000")
port map (
combout => \GRLFPC2_0.N_2888\,
dataf => N_80,
datae => N_70,
datad => \GRLFPC2_0.N_925\,
datac => N_73,
datab => N_69);
GRLFPC2_0_RS1D_CNST_0_A2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000c00000000000")
port map (
combout => \GRLFPC2_0.RS1D_CNST\,
dataf => \GRLFPC2_0.N_2888\,
datae => N_72,
datad => N_71,
datac => N_81,
datab => N_74);
GRLFPC2_0_COMB_RS1D_1_U: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff3ff0c000000")
port map (
combout => \GRLFPC2_0.COMB.RS1D_1\,
dataf => \GRLFPC2_0.RS1D_CNST\,
datae => \GRLFPC2_0.COMB.FPDECODE.RS1D5\,
datad => \GRLFPC2_0.N_884\,
datac => N_80,
datab => N_81);
\GRLFPC2_0_COMB_RS1_1_1_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f00f000000000000")
port map (
combout => \GRLFPC2_0.N_2991\,
dataf => N_77,
datae => \GRLFPC2_0.COMB.FPDECODE.ST\,
datad => N_70,
datac => N_69);
\GRLFPC2_0_COMB_RS1_1_1_RNIOBMO_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfffcf00c0ffc000")
port map (
combout => N_36304,
dataf => \GRLFPC2_0.R.A.RS1\(0),
datae => \GRLFPC2_0.N_2989\,
datad => \GRLFPC2_0.N_889\,
datac => N_9,
datab => N_64);
\GRLFPC2_0_COMB_RS1_1_1_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f00f000000000000")
port map (
combout => \GRLFPC2_0.N_2993\,
dataf => N_79,
datae => \GRLFPC2_0.COMB.FPDECODE.ST\,
datad => N_70,
datac => N_69);
\GRLFPC2_0_COMB_RS1_1_1_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f00f000000000000")
port map (
combout => \GRLFPC2_0.N_2990\,
dataf => N_76,
datae => \GRLFPC2_0.COMB.FPDECODE.ST\,
datad => N_70,
datac => N_69);
\GRLFPC2_0_COMB_RS1_1_1_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f00f000000000000")
port map (
combout => \GRLFPC2_0.N_2992\,
dataf => N_78,
datae => \GRLFPC2_0.COMB.FPDECODE.ST\,
datad => N_70,
datac => N_69);
\GRLFPC2_0_COMB_RS1_1_1_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f00f000000000000")
port map (
combout => \GRLFPC2_0.N_2989\,
dataf => N_75,
datae => \GRLFPC2_0.COMB.FPDECODE.ST\,
datad => N_70,
datac => N_69);
GRLFPC2_0_COMB_RSDECODE_UN1_FPCI_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000f0000")
port map (
combout => \GRLFPC2_0.COMB.RSDECODE.UN1_FPCI_2\,
dataf => N_60,
datae => N_55,
datad => N_63,
datac => N_62);
GRLFPC2_0_COMB_RSDECODE_UN1_FPCI_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ff00")
port map (
combout => \GRLFPC2_0.COMB.RSDECODE.UN1_FPCI_1\,
dataf => N_59,
datae => N_56,
datad => N_61);
GRLFPC2_0_COMB_FPDECODE_RDD6_0_A2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00000000000000")
port map (
combout => \GRLFPC2_0.COMB.FPDECODE.RDD6\,
dataf => \GRLFPC2_0.N_92\,
datae => N_61,
datad => \GRLFPC2_0.N_3418\,
datac => N_56,
datab => N_55);
GRLFPC2_0_RS1V_0_SQMUXA_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffc000000000")
port map (
combout => \GRLFPC2_0.RS1V_0_SQMUXA_1\,
dataf => \GRLFPC2_0.N_620\,
datae => \GRLFPC2_0.N_925\,
datad => \GRLFPC2_0.COMB.FPDECODE.RDD6\,
datac => \GRLFPC2_0.COMB.RSDECODE.UN1_FPCI_2\,
datab => \GRLFPC2_0.COMB.RSDECODE.UN1_FPCI_1\);
GRLFPC2_0_COMB_RS1V_1_IV: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0c0c0c00")
port map (
combout => \GRLFPC2_0.COMB.RS1V_1\,
dataf => \GRLFPC2_0.N_1072_M\,
datae => \GRLFPC2_0.RS1V_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_884\,
datac => N_80,
datab => N_81);
GRLFPC2_0_COMB_RS1V_1_IV_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c300c300c3000000")
port map (
combout => \GRLFPC2_0.N_1072_M\,
dataf => N_83,
datae => N_82,
datad => \GRLFPC2_0.COMB.FPDECODE.ST\,
datac => N_70,
datab => N_69);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_232__G2_0_7612_I_A7_7\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7612_I_A7_7\,
dataf => \GRLFPC2_0.FPCI_O_3\(74),
datae => \GRLFPC2_0.FPCI_O_0\(60),
datad => \GRLFPC2_0.FPCI_O_0\(69),
datac => \GRLFPC2_0.FPCI_O_0\(70));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_232__G2_0_7612_I_A7_10\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0030000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7612_I_A7_10\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7612_I_A7_7\,
datae => \GRLFPC2_0.HOLDN_O\,
datad => \GRLFPC2_0.FPCI_O_0\(59),
datac => \GRLFPC2_0.FPCI_O_0\(63),
datab => \GRLFPC2_0.FPCI_O_0\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_232__G2_0_7612_I_A7_6\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7612_I_A7_6\,
dataf => \GRLFPC2_0.FPCI_O_3\(73),
datae => \GRLFPC2_0.FPCI_O_0\(62),
datad => \GRLFPC2_0.FPCI_O_3\(0),
datac => \GRLFPC2_0.COMB.LOCKGEN.LOCKI_O_3\);
GRLFPC2_0_FPI_LDOP_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffff3000000")
port map (
combout => \GRLFPC2_0.FPI.LDOP_1\,
dataf => \GRLFPC2_0.R.MK.RST\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7612_I_A7_10\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7612_I_A7_6\,
datac => \GRLFPC2_0.R.STATE_O_3\(1),
datab => \GRLFPC2_0.R.STATE_O_3\(0));
\GRLFPC2_0_FPI_OP1_63_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPI.OP1\(63),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => N_630,
datad => N_694);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3639\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_CIN_2_RNIHRRR7: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fccfcffcc00c0cc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_319__G1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_60.Z_1_CO1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1281_I\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_58\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.CIN_2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_SUB_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffff000000ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(19),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(8));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_173_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0c000ccccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(173),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(173));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_14_171_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_14\(171),
dataf => N_59283,
datae => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN7_STKGEN_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3cff3c00c3ffc3")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN7_STKGEN\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10579\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(372),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(371));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIACPP1_314_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3c003c003c003c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5322\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(114),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(372),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(314));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN7_STKGEN_0_RNIE58C2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f300000c0c0c0c")
port map (
combout => N_59285,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.NOTPROP\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN7_STKGEN\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5322\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(373));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_0_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI7UTA_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00f000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_947_I\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(370));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI7UTA_0_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f0ff0fff0f00f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SALSBS_2\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(370));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI3UVA_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0cf3f30cf30cf30c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SALSBS_1\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(369));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00fff0f00000f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(312));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIFSVE_24_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fffff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5446\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10579\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(313));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN2_MIXOIN_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00f0000000f0")
port map (
combout => N_59284,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.GEN\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.NOTPROP\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(373));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN2_MIXOIN_1_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcfff3fffcccc000")
port map (
combout => N_59286,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN13_GEN\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_947_I\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5324\,
datac => N_59284,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SALSBS_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN2_MIXOIN_1_RNI9PST4_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"003c03c03c00c003")
port map (
combout => N_59336,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SBLSBS_1\(1),
datae => N_59286,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_959_I\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SBLSBS_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5452\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNI08K39_315_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0cffffffffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1_2\,
dataf => N_59336,
datae => N_59287,
datad => N_59285,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(315));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_0_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00fff0f00000f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(311));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff00ff000ffff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI3UVA_0_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0c0c000c000c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_1_CO0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(369));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_CIN_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f3cc3f000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6583\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_60_Z_1_CO1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c0ffffc000c0c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_60.Z_1_CO1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_60.Z_1_CO0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_12247\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6583\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2_3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_CIN_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f3cc3f000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5771\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_60_Z_1_CO0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff00ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_60.Z_1_CO0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_2_1_CO1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_CIN_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03fcf30c00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6961\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_CIN_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f33f0cc00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.CIN_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6961\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(57),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(316));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10634\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(258));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_12_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3330303033000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2267\,
dataf => N_33001_1,
datae => N_33133_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2485\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2538\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0003000c0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2351\,
dataf => N_32032_I,
datae => N_31921_1_0,
datad => N_32203_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2525\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_0_A2_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3f0033000f000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8752\,
dataf => N_32032_I,
datae => N_31725_1_0,
datad => N_32120_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_O2_1_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00030000c0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_339\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_O2_39_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffcf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_523\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2405\,
datae => N_31725_1_0,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2490\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2518\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2546\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_0_O2_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf0cc00f0f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8695\,
dataf => N_33133_1,
datae => N_32619_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2508\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2536\,
datab => N_32434_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_62_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffc0c0c0ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_568\,
dataf => N_32340_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2513\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2490\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2485\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2484\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_2_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cccc0c00cccc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2671\,
dataf => N_31886_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2504\,
datad => N_31924_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_O2_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffcccfffff000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_726\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2779\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2534\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_20_0\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2484\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_X3_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_885_I\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\(78));
GRLFPC2_0_COMB_UN1_R_A_RS1_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0c0c0c0c0c0c0c")
port map (
combout => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
dataf => \GRLFPC2_0.N_27\,
datae => \GRLFPC2_0.N_7\,
datad => \GRLFPC2_0.COMB.UN1_FPCI_3_1\,
datac => \GRLFPC2_0.R.A.RS1D\,
datab => \GRLFPC2_0.R.A.RS1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_PCTRL_1_SUM_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ffff00ffff0000")
port map (
combout => N_28947,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_PCTRL_1_SUM_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3fc0ff00ff00ff00")
port map (
combout => N_28952,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_1_2_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000000000000")
port map (
combout => N_27776_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_27_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff0000000000")
port map (
combout => N_31743,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O18_2_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0000ff000000ff")
port map (
combout => N_31703,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O18_3_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00000000ffff00")
port map (
combout => N_31704,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O9_0_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff000000")
port map (
combout => N_31753,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O13_7_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00300c03000000")
port map (
combout => N_31803,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_X2_58_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffff0000")
port map (
combout => N_32022_I,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_16_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00000000ff0000")
port map (
combout => N_32232,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_X2_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffff0000")
port map (
combout => N_32885_I,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_4_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_32230,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_5_0_12_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_32052_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_X2_1_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffff0000")
port map (
combout => N_28030_I,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_33071_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_X2_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffff0000")
port map (
combout => N_32662_I,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A2_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_31921_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A28_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c00000cc00000000")
port map (
combout => N_33055,
dataf => N_31921_1,
datae => N_31766_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_X4_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffff0000")
port map (
combout => N_33043_I,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O17_4_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030000cc0c00f00")
port map (
combout => N_33193,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_32141_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_1_1_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9074_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84));
GRLFPC2_0_COMB_V_MK_BUSY_2_4: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000f0000000000")
port map (
combout => \GRLFPC2_0.R.MK.BUSY_4\,
dataf => \GRLFPC2_0.FPO.BUSY_O_0\,
datae => \GRLFPC2_0.R.MK.RST2_O_0\,
datad => \GRLFPC2_0.R.MK.HOLDN1_O_0\,
datac => \GRLFPC2_0.COMB.ANNULFPU_1_O_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A2_1_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_32425_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_1_1_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_31725_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_8_1_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_33063_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_1_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f00cc0000000000")
port map (
combout => N_31864,
dataf => N_31921_1_0,
datae => N_31774_1,
datad => N_31864_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_2_2_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_31767_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_X2_0_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffff0000")
port map (
combout => N_32390_I,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_15_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_31865_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_X2_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffff0000")
port map (
combout => N_31691_I,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_19_1_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_31940_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A20_1_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_32140_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A20_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330c000000000000")
port map (
combout => N_32483,
dataf => N_32032_I,
datae => N_33372,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_I_0_O26_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000ffff")
port map (
combout => N_32020,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_9_1_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_32131_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A28_1_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_31718_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_3_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c0cf000000000000")
port map (
combout => N_32904,
dataf => N_32932,
datae => N_31941_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_7_1_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_31886_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_7_1_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_28591_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_11_1_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_33076_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A2_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_32705_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_0_1_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_32645_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_3_1_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_32343_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_5_2_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_32050_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_0_1_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_32047_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A17_1_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_32550_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_31769_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_4_1_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_32708_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_5_1_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_32620_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_6_2_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_32422_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_10_1_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_32435_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_13_1_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_31919_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A12_1_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_31715_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_1_1_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_32632_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_1_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000330000000000")
port map (
combout => N_33312,
dataf => N_32632_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(81),
datad => N_33312_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_2_1_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_27929_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_9_1_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_31989_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_6_1_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_31819_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_3_1_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_33136_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_3_2_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00ff00ff")
port map (
combout => N_31718_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_8_1_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_27297_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_O2_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000ffff")
port map (
combout => N_33232,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A24_1_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_32015_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_23_1_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_33057_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_31768_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A15_1_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_31808_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_3_2_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_32340_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_7_1_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_32438_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_MIFROMINST_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00f00033003300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.MIFROMINST_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(73),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(71),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(74));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_26_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30f0303000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2722\,
dataf => N_32032_I,
datae => N_31725_1_0,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_320\,
datac => N_32120_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000c00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW_6\(0),
dataf => N_61,
datae => N_59,
datad => N_62,
datac => N_58,
datab => N_57);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_X2_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffff0000")
port map (
combout => N_27758_I,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_1_1_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_31864_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_X2_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffff0000")
port map (
combout => N_31899_I,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_22_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_22__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_1_2\(22),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1071\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2640\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_20_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffff0f000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_20__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1931\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2763\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2485\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2484\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_1_1_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_31819_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_2_1_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_32136_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_1_RNIBC2F_9_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcccf000cccc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19\(9),
dataf => N_33001_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1967_1\,
datad => N_32434_2,
datac => N_31924_1,
datab => N_32136_1);
GRLFPC2_0_COMB_FPDECODE_FPOP3_0_A2_0_RNIDE201_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000c000000")
port map (
combout => \GRLFPC2_0.R.A.LD_0_0_G1_0\,
dataf => N_71,
datae => \GRLFPC2_0.N_77\,
datad => N_81,
datac => N_73,
datab => N_80);
GRLFPC2_0_COMB_RDD_1_M14_0_A2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00000000000000")
port map (
combout => \GRLFPC2_0.N_73\,
dataf => \GRLFPC2_0.R.A.LD_0_0_G1_0\,
datae => N_70,
datad => N_69);
GRLFPC2_0_COMB_RDD_1_M14_0_A2_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000c000000")
port map (
combout => \GRLFPC2_0.N_78\,
dataf => N_57,
datae => N_58,
datad => \GRLFPC2_0.N_37\,
datac => N_56,
datab => N_61);
GRLFPC2_0_COMB_RDD_1_M14_0_O2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00000c00")
port map (
combout => \GRLFPC2_0.N_40\,
dataf => \GRLFPC2_0.N_78\,
datae => N_62,
datad => \GRLFPC2_0.N_38\,
datac => N_55,
datab => N_56);
GRLFPC2_0_R_X_AFSR_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f00000000")
port map (
combout => \GRLFPC2_0.R.X.AFSR_0_0_G1\,
dataf => \GRLFPC2_0.R.E.AFSR_O\,
datae => \GRLFPC2_0.N_1829_O\,
datad => N_291,
datac => N_292);
GRLFPC2_0_R_X_AFQ_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f00000000")
port map (
combout => \GRLFPC2_0.R.X.AFQ_0_0_G1\,
dataf => \GRLFPC2_0.R.E.AFQ_O\,
datae => \GRLFPC2_0.N_1829_O\,
datad => N_291,
datac => N_292);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_13_1_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_32627_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_5_1_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_32688_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_3_1_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_32786_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_1_1_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_32124_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_M20_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => N_32327,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A22_1_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_32064_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A12_1_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_32645_3,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_11_1_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_31999_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_X2_1_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffff0000")
port map (
combout => N_32032_I,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O2_3_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0f0000cccc00cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_377\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(76),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(71),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(74));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A2_5_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f033ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2457\,
dataf => N_28949,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(71),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(74));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_X2_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffff0000")
port map (
combout => N_32530_I,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_5_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c0c00000f0c03000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_5\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_255\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2494\,
datad => N_32487_2,
datac => N_32530_I,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_2_1_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_32272_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_9_1_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_31775_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84));
GRLFPC2_0_COMB_RDD_1_M14_0_O2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffff0000")
port map (
combout => \GRLFPC2_0.N_37\,
dataf => N_60,
datae => N_62,
datad => N_55);
GRLFPC2_0_COMB_V_MK_RST_1_4: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000f00000")
port map (
combout => \GRLFPC2_0.R.MK.RST_4\,
dataf => \GRLFPC2_0.R.MK.RST2\,
datae => \GRLFPC2_0.R.MK.HOLDN2\,
datad => \GRLFPC2_0.R.MK.RST2_O\,
datac => \GRLFPC2_0.COMB.ANNULFPU_1_O\);
GRLFPC2_0_COMB_V_MK_RST_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000000000000000")
port map (
combout => \GRLFPC2_0.R.MK.RST\,
dataf => \GRLFPC2_0.FPO.BUSY_O\,
datae => \GRLFPC2_0.R.MK.RST_4\,
datad => \GRLFPC2_0.HOLDN_O\,
datac => \GRLFPC2_0.R.MK.HOLDN2_O\);
GRLFPC2_0_FPI_START: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000f000000000")
port map (
combout => \GRLFPC2_0.FPI.START\,
dataf => \GRLFPC2_0.N_1000\,
datae => \GRLFPC2_0.R.MK.RST\,
datad => \GRLFPC2_0.R.MK.RST2\,
datac => N_9);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MAPMULXFF_UN7_UNIMPMAP_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ffffff0f000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MAPMULXFF.UN7_UNIMPMAP\,
dataf => N_69,
datae => N_61,
datad => N_59,
datac => N_62);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_ENA_67_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"030303030303ff00")
port map (
combout => N_48774,
dataf => \GRLFPC2_0.FPI.START\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(67),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MAPMULXFF.UN7_UNIMPMAP\,
datab => N_63);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNI654D_67_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2645\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(67));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_RESULT_IV_RNO_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000c30000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SFTLFT.AREGXORBREG_I_M\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_27_S_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(12),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(13));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_A3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccc0c0cc00c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2477\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_318\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422\,
datad => N_31813_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(66));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A21_1_59_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_31762_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O2_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00cc00ff0fcc0c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O2_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_647\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_A3_0_1\,
datac => N_32136_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffcccf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2477\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O2_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2765\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_13_1_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_31996_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_11_1_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_32136_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_PCTRL_1_CO2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0f0000000f000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2757\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(71),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(74),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(63));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_O3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0000033330033")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_329\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(76),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(71),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(74));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_O28_5_60_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000ffff")
port map (
combout => N_33040,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_1_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_31838_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_6_1_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_32120_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_9_1_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_32775_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_32434_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_6_3_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffff3ffffff33")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_6_3\(4),
dataf => N_31921_1_0,
datae => N_32141_1_0,
datad => N_32775_1,
datac => N_32434_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(67));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_3_0_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_31924_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(78));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_51_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0f0f0f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2555\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_318\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O2_2\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O2_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(66));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_UN10_SELECTEDMIPTR_I_0_O2_RNI5AT05: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000c00c00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3729_I_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5088\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2807\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNI21Q11_76_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_237\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(76));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_27_S_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_27_S_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(49),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(51));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_24: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"66666666e6e6e666")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10927\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV\,
datae => \GRLFPC2_0.FPO.FRAC\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN30_CONDITIONAL_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(48));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_21: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f00f0f0ff0f00ff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10924\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI0TK9GF3_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2\,
dataf => N_26592,
datae => N_26591,
datad => N_26534);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_10: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0000fff00ff00f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10913\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(12),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_6: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f03cc30f0f3cc3")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10909\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\(12),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(13));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0000ff00ff00ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10906\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(48));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_15: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbea7362d9c85140")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10918\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10909\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10916\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10906\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10913\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIP28I_252_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4167_I_0_I_A3_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(256),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(254),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(255),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(252));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIC5G41_250_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000300000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4167_I_0_I_A3_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4167_I_0_I_A3_4\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(251),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(257),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(250),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(253));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIC36J3_246_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffcfffccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2807\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1919\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4167_I_0_I_A3_6\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_529\,
datac => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_46_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(46),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_45_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(45),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_40_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(40),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_39_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(39),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_38_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(38),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_37_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(37),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_36_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(36),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_50: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"1428000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_50\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_42\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_27\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(30),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(30),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(47),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_35_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(35),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_44_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(44),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_41_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(41),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(55),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(51),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(50),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_49: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0660000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_49\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_40\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_23\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(47),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(35));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_49_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(49),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(48),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(57),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f00f0fcc0033ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(57),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(174));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(56),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_42_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(42),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(52),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_32_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(32),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_28_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff000f0ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(28),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_20_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff000f0ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(20),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff000f0ffc000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_14: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f00f00f00f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_14\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(15),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_36: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03000c003000c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_36\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(28),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(20),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_14\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(20));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f00f00f00f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(16),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(16));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_53: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"6000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_53\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_38\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_36\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_39\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_19_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0ff00f0f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(19),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_12: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f00f00f00f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_12\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(10),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff000f0ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(27),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_26_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff000f0ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(26),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_10: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f00f00f00f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_10\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(26),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_23_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff000f0ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(23),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_22_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0ff00f0f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(22),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_21_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff000f0ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(21),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_4: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f0f0000f0f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(21),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(21));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_31: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"030c30c000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_31\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_4\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(23),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(22),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(23),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(54),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_52: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"1428000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_52\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_46\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_31\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff000f0ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(25),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_24_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff000f0ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(24),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_8: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f0f0000f0f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(8));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_6: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f00f00f00f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_32: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"030c30c000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_32\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_45: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"1020408000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_45\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_32\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(24),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_8\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(34),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(33),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff000f0ffc000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(114),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff000f0ffc000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(115),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0003030000303000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5410\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5391\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_37: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000012480000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_37\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN18_XZXBUS_14\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(33));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"8000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_52\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_53\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_50\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_49\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_45\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_37\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI85QEL01_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_176__G2\,
dataf => N_26534,
datae => N_26588,
datad => N_26587);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI4DONJ53_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_175__G2\,
dataf => N_26534,
datae => N_26590,
datad => N_26589);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10879\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(243),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(256));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_1_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10866\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10878\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(257));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_9_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff03cf0f0f03cf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(9),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(9),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_9_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10887\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(248));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff03cf0f0f03cf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(9),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(237));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_7_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10885\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(237),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(250));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff03cf0f0f03cf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(238));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10884\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(238),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(251));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10883\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(239),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(252));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5339\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(232));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_12_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10890\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(232),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(245));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5301\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_10_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10888\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(247));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5343\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_11_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10889\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff0f0f03cf03cf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(240));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10882\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(240),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(253));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_1_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10869\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff03cf0f0f03cf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(8),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(9),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10886\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(249));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPYBUS_2_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_5: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff9")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_8\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10881\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(241),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(254));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPYBUS_2_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ffffff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_8: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffd827")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_6\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10868\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10881\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10880\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(255));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_1_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10867\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_NE: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffd827")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_I\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_10\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_8\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10867\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10880\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN30_CONDITIONAL_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN30_CONDITIONAL_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5330\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\(12),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_I\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIC1BA6U1_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(54),
dataf => N_26534,
datae => N_26586,
datad => N_26585);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIKMVUAK2_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(52),
dataf => N_26534,
datae => N_26582,
datad => N_26581);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIGF3OUC2_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(53),
dataf => N_26534,
datae => N_26584,
datad => N_26583);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI4S44SP_50_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(50),
dataf => N_26534,
datae => N_26578,
datad => N_26577);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI8QD21O2_51_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(51),
dataf => N_26534,
datae => N_26580,
datad => N_26579);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNICDLPFJ2_47_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(47),
dataf => N_26534,
datae => N_26572,
datad => N_26571);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI4D0LPQ1_49_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(49),
dataf => N_26534,
datae => N_26576,
datad => N_26575);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI8DED8B2_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(48),
dataf => N_26534,
datae => N_26574,
datad => N_26573);
GRLFPC2_0_COMB_FPDECODE_RDD6_0_A2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff0000000000")
port map (
combout => \GRLFPC2_0.N_92\,
dataf => N_60,
datae => N_57,
datad => N_58);
GRLFPC2_0_COMB_FPDECODE_RDD5_0_A2_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000ff")
port map (
combout => \GRLFPC2_0.N_3418\,
dataf => N_59,
datae => N_63,
datad => N_62);
GRLFPC2_0_UN1_MOV_1_SQMUXA_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff000c00ff000000")
port map (
combout => \GRLFPC2_0.UN1_MOV_1_SQMUXA_0\,
dataf => \GRLFPC2_0.MOV_2_SQMUXA_1\,
datae => \GRLFPC2_0.N_925\,
datad => \GRLFPC2_0.N_620\,
datac => N_55,
datab => N_56);
GRLFPC2_0_UN1_MOV_1_SQMUXA_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => \GRLFPC2_0.N_909_7\,
dataf => \GRLFPC2_0.N_93\,
datae => N_62,
datad => N_57,
datac => N_58,
datab => N_59);
GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_7_4: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000f")
port map (
combout => \GRLFPC2_0.COMB.FPDECODE.UN1_FPCI_7_4\,
dataf => N_60,
datae => N_55,
datad => N_59,
datac => N_58);
GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_7: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000000000000000")
port map (
combout => \GRLFPC2_0.N_908_7\,
dataf => \GRLFPC2_0.COMB.FPDECODE.UN1_FPCI_7_4\,
datae => N_62,
datad => N_61,
datac => N_57,
datab => N_56);
GRLFPC2_0_UN1_MOV_1_SQMUXA: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000fc00")
port map (
combout => \GRLFPC2_0.N_896\,
dataf => \GRLFPC2_0.UN1_MOV_1_SQMUXA_0\,
datae => N_63,
datad => \GRLFPC2_0.N_620\,
datac => \GRLFPC2_0.N_909_7\,
datab => \GRLFPC2_0.N_908_7\);
GRLFPC2_0_COMB_PEXC8_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => CPO_EXCZ,
dataf => \GRLFPC2_0.R.STATE\(0),
datae => \GRLFPC2_0.R.STATE\(1));
GRLFPC2_0_COMB_LOCKGEN_LOCKI_I_0_RNIHL981: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff000000")
port map (
combout => \GRLFPC2_0.N_1000\,
dataf => \GRLFPC2_0.COMB.LOCKGEN.LOCKI_I_I\,
datae => \GRLFPC2_0.N_939_I_0_A2_2\,
datad => \GRLFPC2_0.N_889\);
GRLFPC2_0_COMB_UN1_FPCI_3_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00000000000000")
port map (
combout => \GRLFPC2_0.COMB.UN1_FPCI_3_1\,
dataf => \GRLFPC2_0.COMB.FPDECODE.ST_O\,
datae => \GRLFPC2_0.R.A.RS1D\,
datad => N_152);
GRLFPC2_0_COMB_UN1_FPCI_3_1_0_O2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000ffff")
port map (
combout => \GRLFPC2_0.N_7\,
dataf => \GRLFPC2_0.R.STATE_O\(1),
datae => \GRLFPC2_0.R.STATE_O\(0));
GRLFPC2_0_R_A_AFQ_RET_2_RNIMUGP: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000f")
port map (
combout => \GRLFPC2_0.N_27\,
dataf => \GRLFPC2_0.FPCI_O\(74),
datae => \GRLFPC2_0.FPCI_O\(73),
datad => \GRLFPC2_0.FPCI_O\(0),
datac => \GRLFPC2_0.COMB.LOCKGEN.LOCKI_O\);
GRLFPC2_0_COMB_UN1_FPCI_4: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0c0c0c0c0c0c0c")
port map (
combout => \GRLFPC2_0.COMB.UN1_FPCI_4\,
dataf => \GRLFPC2_0.N_27\,
datae => \GRLFPC2_0.N_7\,
datad => \GRLFPC2_0.COMB.UN1_FPCI_3_1\,
datac => \GRLFPC2_0.R.A.RS2D\,
datab => \GRLFPC2_0.R.A.RS2\(0));
GRLFPC2_0_COMB_FPDECODE_RDD5_0_A2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000f00000")
port map (
combout => \GRLFPC2_0.N_93\,
dataf => N_55,
datae => N_56,
datad => N_60,
datac => N_61);
GRLFPC2_0_COMB_FPDECODE_RS1D5_0_A2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000c00")
port map (
combout => \GRLFPC2_0.COMB.FPDECODE.RS1D5\,
dataf => N_63,
datae => N_62,
datad => \GRLFPC2_0.N_93\,
datac => N_58,
datab => N_59);
GRLFPC2_0_COMB_FPDECODE_FPOP3_0_A2_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff0000000000")
port map (
combout => \GRLFPC2_0.N_94\,
dataf => N_73,
datae => N_70,
datad => N_71);
GRLFPC2_0_COMB_LOCKGEN_LOCKI_I_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0300")
port map (
combout => \GRLFPC2_0.COMB.LOCKGEN.LOCKI_I_I\,
dataf => \GRLFPC2_0.COMB.LOCKGEN.LOCKI_I_1\,
datae => \GRLFPC2_0.N_1092\,
datad => \GRLFPC2_0.COMB.SEQERR.UN13_OP_0_3\,
datac => N_73,
datab => N_71);
GRLFPC2_0_COMB_LOCKGEN_UN8_DEPCHECK: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff0")
port map (
combout => \GRLFPC2_0.N_1093\,
dataf => \GRLFPC2_0.R.X.LD\,
datae => \GRLFPC2_0.R.M.LD\,
datad => \GRLFPC2_0.R.A.LD\,
datac => \GRLFPC2_0.R.E.LD\);
GRLFPC2_0_COMB_LOCKGEN_LOCKI_I_0_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3fffffff0fff0")
port map (
combout => \GRLFPC2_0.COMB.LOCKGEN.LOCKI_I_1\,
dataf => \GRLFPC2_0.N_178\,
datae => \GRLFPC2_0.N_1093\,
datad => N_83,
datac => N_82,
datab => \GRLFPC2_0.N_1092\);
GRLFPC2_0_COMB_FPDECODE_FPOP3_0_A2_0_RNIDE201: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00000000000000")
port map (
combout => \GRLFPC2_0.COMB.FPDECODE.ST\,
dataf => N_71,
datae => \GRLFPC2_0.N_77\,
datad => N_81,
datac => N_73,
datab => N_80);
GRLFPC2_0_RS2_0_SQMUXA_0_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff0000000000")
port map (
combout => \GRLFPC2_0.N_889_1\,
dataf => N_74,
datae => N_70,
datad => N_71);
GRLFPC2_0_RS2_0_SQMUXA_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000c0000000000")
port map (
combout => \GRLFPC2_0.N_889\,
dataf => \GRLFPC2_0.N_889_1\,
datae => N_72,
datad => N_73,
datac => N_80,
datab => N_81);
GRLFPC2_0_RS2_0_SQMUXA_0_RNITQP41: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0000")
port map (
combout => \GRLFPC2_0.N_1092\,
dataf => \GRLFPC2_0.N_889\,
datae => \GRLFPC2_0.COMB.FPDECODE.ST\);
GRLFPC2_0_COMB_FPDECODE_FPOP3_0_A2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => \GRLFPC2_0.N_77\,
dataf => N_74,
datae => N_72);
GRLFPC2_0_COMB_SEQERR_UN13_OP_0_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cf00000000000000")
port map (
combout => \GRLFPC2_0.COMB.SEQERR.UN13_OP_0_3\,
dataf => \GRLFPC2_0.N_77\,
datae => N_81,
datad => N_80,
datac => N_70,
datab => N_69);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_6_1_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_27553_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_6_1_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_31724_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_6_1_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_32069_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_4_2_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000000000000")
port map (
combout => N_32841_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_3_1_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_31774_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_7_2_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_32712_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_4_1_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_32566_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A20_1_48_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_31765_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_0_1_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_32220_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_7_2_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_31723_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A29_1_57_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_31941_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_13_2_34_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_28580_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_4_2_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_31813_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_3_1_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_32070_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_8_1_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_32487_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_14_1_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_31766_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_O2_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffffffff")
port map (
combout => N_33298,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A2_33_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_32066_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_0_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffffffff")
port map (
combout => N_33176,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O24_0_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0000")
port map (
combout => N_32739,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A2_55_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_31839_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_I_O2_31_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffffffff")
port map (
combout => N_31892,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_X2_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffff0000")
port map (
combout => N_32673_I,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O22_2_53_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_320\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_15_1_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_32203_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A25_1_54_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_32908_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_13_2_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_31766_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_X2_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffff0000")
port map (
combout => N_32394_I,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_9_1_52_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_33136_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_O28_16_56_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00000000ff00ff")
port map (
combout => N_32405,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A2_13_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_31763_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_6_1_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_32142_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_O2_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_247\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_0_1_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_32048_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_6_1_18_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_33138_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O13_1_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000ffff")
port map (
combout => N_31788,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_O2_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000ffff")
port map (
combout => N_31688,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNI5MLD_247_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_529\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(248),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(249),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(247));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIP28I_0_252_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_I_0_A2_4\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(256),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(254),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(255),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(252));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_OPREXCSHFT_UN14_EXMIPTRLSBS: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000030300ff03ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN14_EXMIPTRLSBS\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_6\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1919\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3848\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2726\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN26_NOTAINFNAN_4: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN26_NOTAINFNAN_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(238),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(241),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(239),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(240));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN26_NOTAINFNAN_RNIS40K: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000f0f0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5065\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7144\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3848\,
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNI8E7I_239_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_4\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(243),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(241),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(239));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIHOE41_237_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_6\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_4\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(238),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(237),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(240));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN3_NOTAZERODENORM: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3848\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_1_RNI09QD1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000c0000000")
port map (
combout => N_81626,
dataf => N_81619,
datae => \GRLFPC2_0.FPO.EXP\(4),
datad => \GRLFPC2_0.FPO.EXP\(1),
datac => \GRLFPC2_0.FPO.EXP\(3),
datab => \GRLFPC2_0.FPO.EXP\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0cccc0f00cccc")
port map (
combout => N_80628,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10080\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10140\,
datac => N_76344,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_12_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0cccc0f00cccc")
port map (
combout => N_80616,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10070\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10130\,
datac => N_76344,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN1_CCIN_RNI0OHDB: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c00000c0003f3f00")
port map (
combout => N_81684,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SCLSBS_2\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SCLSBS_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_954\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7210\);
N_81985 <= not N_56;
N_81986 <= not \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datain => N_80674,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_9_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datain => N_80673,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_18_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18),
datain => N_80672,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_19_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19),
datain => N_80671,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_20_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datain => N_80670,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_21_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
datain => N_80669,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_22_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22),
datain => N_80668,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_23_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datain => N_80667,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_24_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24),
datain => N_80666,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_25_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datain => N_80665,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_26_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26),
datain => N_80664,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_27_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27),
datain => N_80663,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_28_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28),
datain => N_80662,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_29_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29),
datain => N_80661,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_30_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30),
datain => N_80660,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_31_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31),
datain => N_80659,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_32_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32),
datain => N_80658,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_33_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33),
datain => N_80657,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_34_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34),
datain => N_80656,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_35_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datain => N_80655,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_36_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36),
datain => N_80654,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_37_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37),
datain => N_80653,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_38_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
datain => N_80652,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_39_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39),
datain => N_80651,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_40_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
datain => N_80650,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_41_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41),
datain => N_80649,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_42_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42),
datain => N_80648,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_43_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43),
datain => N_80647,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_44_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44),
datain => N_80646,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_45_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45),
datain => N_80645,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_46_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46),
datain => N_80644,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_47_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47),
datain => N_80643,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_48_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48),
datain => N_80642,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_49_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
datain => N_80641,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_50_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datain => N_80640,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_51_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datain => N_80639,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_52_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datain => N_80638,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_53_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datain => N_80637,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_54_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datain => N_80636,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_55_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datain => N_80635,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_56_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
datain => N_80634,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_57_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datain => N_80633,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_3_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datain => N_80632,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_0: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7782_1\,
datain => N_80631,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_10_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
datain => N_80630,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_16_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16),
datain => N_80629,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_2_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datain => N_80628,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_13_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13),
datain => N_80627,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_4_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4),
datain => N_80626,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_6_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6),
datain => N_80625,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_2: stratixii_lcell_ff port map (
regout => N_79982,
datain => N_80624,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_15_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
datain => N_80623,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_5_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
datain => N_80622,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_11_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11),
datain => N_80621,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_17_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datain => N_80620,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_11: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_10\,
datain => N_80619,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_7_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7),
datain => N_80618,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_8_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
datain => N_80617,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_12_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12),
datain => N_80616,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_14_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14),
datain => N_80615,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_20: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_9\,
datain => N_80614,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_122: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(101),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(101),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_113: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(100),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(100),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_110: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(77),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(77),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_104: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(99),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(99),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_112_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(112),
clk => N_8,
sload => \GRLFPC2_0.FPI.LDOP_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(112),
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	ena => VCC);
\GRLFPC2_0.FPI.LDOP_I\ <= not \GRLFPC2_0.FPI.LDOP_4\;
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_111_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(111),
clk => N_8,
sload => \GRLFPC2_0.FPI.LDOP_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(111),
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_110_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(110),
clk => N_8,
sload => \GRLFPC2_0.FPI.LDOP_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(110),
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_109_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(109),
clk => N_8,
sload => \GRLFPC2_0.FPI.LDOP_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(109),
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_108_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(108),
clk => N_8,
sload => \GRLFPC2_0.FPI.LDOP_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(108),
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_107_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(107),
clk => N_8,
sload => \GRLFPC2_0.FPI.LDOP_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(107),
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_82_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(82),
clk => N_8,
sload => \GRLFPC2_0.FPI.LDOP_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(82),
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_83_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(83),
clk => N_8,
sload => \GRLFPC2_0.FPI.LDOP_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(83),
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_102_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(102),
clk => N_8,
sload => \GRLFPC2_0.FPI.LDOP_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(102),
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_79_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(79),
clk => N_8,
sload => \GRLFPC2_0.FPI.LDOP_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(79),
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_78_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(78),
clk => N_8,
sload => \GRLFPC2_0.FPI.LDOP_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(78),
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_73_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(73),
clk => N_8,
sload => \GRLFPC2_0.FPI.LDOP_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(73),
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_75_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(75),
clk => N_8,
sload => \GRLFPC2_0.FPI.LDOP_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(75),
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_96_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(96),
clk => N_8,
sload => \GRLFPC2_0.FPI.LDOP_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(96),
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_93_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(93),
clk => N_8,
sload => \GRLFPC2_0.FPI.LDOP_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(93),
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_69_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(69),
clk => N_8,
sload => \GRLFPC2_0.FPI.LDOP_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(69),
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_71_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(71),
clk => N_8,
sload => \GRLFPC2_0.FPI.LDOP_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(71),
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_70_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(70),
clk => N_8,
sload => \GRLFPC2_0.FPI.LDOP_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(70),
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_67_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(67),
clk => N_8,
sload => \GRLFPC2_0.FPI.LDOP_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(67),
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_66_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(66),
clk => N_8,
sload => \GRLFPC2_0.FPI.LDOP_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(66),
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_65_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(65),
clk => N_8,
sload => \GRLFPC2_0.FPI.LDOP_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(65),
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_61_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(61),
clk => N_8,
sload => \GRLFPC2_0.FPI.LDOP_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(61),
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_63_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(63),
clk => N_8,
sload => \GRLFPC2_0.FPI.LDOP_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(63),
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_64_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(64),
clk => N_8,
sload => \GRLFPC2_0.FPI.LDOP_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(64),
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_62_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(62),
clk => N_8,
sload => \GRLFPC2_0.FPI.LDOP_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(62),
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_129: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(73),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(73),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_128: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_4_0_RETO\(4),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_4_0\(4),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_127: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2462_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2462\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_251: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(40),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_250: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(98),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_249: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPO.FRAC_RETO\(15),
datain => \GRLFPC2_0.FPO.FRAC\(15),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_248: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPO.FRAC_RETO\(17),
datain => \GRLFPC2_0.FPO.FRAC\(17),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_245: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(39),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_244: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(97),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_243: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPO.FRAC_RETO\(16),
datain => \GRLFPC2_0.FPO.FRAC\(16),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_239: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(18),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_238: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(76),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_237: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPO.FRAC_RETO\(37),
datain => \GRLFPC2_0.FPO.FRAC\(37),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_233: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(37),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_232: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(95),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_231: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPO.FRAC_RETO\(18),
datain => \GRLFPC2_0.FPO.FRAC\(18),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_230: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPO.FRAC_RETO\(20),
datain => \GRLFPC2_0.FPO.FRAC\(20),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_227: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(16),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_226: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(74),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_225: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPO.FRAC_RETO\(41),
datain => \GRLFPC2_0.FPO.FRAC\(41),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_224: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPO.FRAC_RETO\(39),
datain => \GRLFPC2_0.FPO.FRAC\(39),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_221: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(36),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_220: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(94),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_219: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPO.FRAC_RETO\(19),
datain => \GRLFPC2_0.FPO.FRAC\(19),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_218: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPO.FRAC_RETO\(21),
datain => \GRLFPC2_0.FPO.FRAC\(21),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_215: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(34),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_214: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(92),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_212: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPO.FRAC_RETO\(23),
datain => \GRLFPC2_0.FPO.FRAC\(23),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_209: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(33),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_208: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(91),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_207: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPO.FRAC_RETO\(22),
datain => \GRLFPC2_0.FPO.FRAC\(22),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_206: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPO.FRAC_RETO\(24),
datain => \GRLFPC2_0.FPO.FRAC\(24),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_203: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(10),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_202: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(68),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_201: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPO.FRAC_RETO\(45),
datain => \GRLFPC2_0.FPO.FRAC\(45),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_200: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPO.FRAC_RETO\(47),
datain => \GRLFPC2_0.FPO.FRAC\(47),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_198: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_197: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(32),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_196: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(90),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_194: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPO.FRAC_RETO\(25),
datain => \GRLFPC2_0.FPO.FRAC\(25),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_193: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_191: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(31),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_190: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(89),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_188: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPO.FRAC_RETO\(26),
datain => \GRLFPC2_0.FPO.FRAC\(26),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_185: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(30),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_184: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(88),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_182: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPO.FRAC_RETO\(27),
datain => \GRLFPC2_0.FPO.FRAC\(27),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_179: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(29),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_178: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(87),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_176: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPO.FRAC_RETO\(28),
datain => \GRLFPC2_0.FPO.FRAC\(28),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_173: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(60),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_172: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(2),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_171: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_176__G2_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_176__G2\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_170: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPO.FRAC_RETO\(53),
datain => \GRLFPC2_0.FPO.FRAC\(53),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_167: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(59),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_166: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(1),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_165: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_175__G2_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_175__G2\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_164: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPO.FRAC_RETO\(54),
datain => \GRLFPC2_0.FPO.FRAC\(54),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_161: stratixii_lcell_ff port map (
regout => N_26563_RETO,
datain => N_26563,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_160: stratixii_lcell_ff port map (
regout => N_26564_RETO,
datain => N_26564,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_158: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(72),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_156: stratixii_lcell_ff port map (
regout => N_26559_RETO,
datain => N_26559,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_155: stratixii_lcell_ff port map (
regout => N_26560_RETO,
datain => N_26560,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_154: stratixii_lcell_ff port map (
regout => N_26534_RETO,
datain => N_26534,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_153: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(14),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_126: stratixii_lcell_ff port map (
regout => N_55054_RETO,
datain => N_55054,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_125: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_124: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(50),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(50),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_123: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10918_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10918\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_122: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_27_S_0_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_27_S_0\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_121: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(49),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(49),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_120: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10927_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10927\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_118: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_2: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2466_1_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2466_1\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_113: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_112: stratixii_lcell_ff port map (
regout => N_28949_RETO,
datain => N_28949,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_111: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(4),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT\(4),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_110: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_109: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_105: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO(6),
datain => N_56,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_104: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_377_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_377\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_103: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_13_C_RETO\(4),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_13_C\(4),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_98: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_I_0_0_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_I_0_0\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_97: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5330_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5330\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_96: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_RETO\(12),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\(12),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_30: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_1: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(60),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(60),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_54: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0_RETO\(9),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0\(9),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_26: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(58),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(58),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_91: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1164_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1164\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_20: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2474_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2474\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_89: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_237_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_237\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_88: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(77),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_87: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_13: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G1_1\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G1_1_RETI\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_374_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(374),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(374),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_15_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(15),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(15),
clk => N_8,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(9),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(9),
clk => N_8,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_231_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(231),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(231),
clk => N_8,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(11),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(11),
clk => N_8,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(12),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(12),
clk => N_8,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_22: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_RETO\(1),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV\(1),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_79: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(55),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_38: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(54),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_78: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(53),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_151: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(85),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(85),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_149: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(85),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(85),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_148: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(86),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(86),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_146: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(86),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(86),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_145: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(84),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(84),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_143: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(84),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(84),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_142: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(106),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(106),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_140: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(106),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(106),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_139: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(105),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(105),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_137: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(105),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(105),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_136: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(104),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(104),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_135: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_134: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(104),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(104),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_133: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(81),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(81),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_131: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(81),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(81),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_130: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(103),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(103),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_128: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(103),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(103),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_127: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(80),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(80),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_125: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(80),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(80),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_124: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(101),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(101),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_121: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPI.LDOP_RETO\,
datain => \GRLFPC2_0.FPI.LDOP_4\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_120: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(84),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(84),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_117: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(85),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(85),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_115: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(100),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(100),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_112: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(77),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(77),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_108: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(86),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(86),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_106: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(99),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(99),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_103: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(98),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(98),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_99: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(97),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(97),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_97: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(76),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(76),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_95: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(106),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(106),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_92: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(81),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(81),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_90: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(95),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(95),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_88: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(74),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(74),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_86: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(105),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(105),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_84: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(80),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(80),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_82: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(94),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(94),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_80: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(104),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(104),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_78: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(103),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(103),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_76: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(101),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(101),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_74: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(89),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(89),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_72: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(88),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(88),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_70: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(92),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(92),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_68: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(77),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(77),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_65: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(91),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(91),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_63: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(68),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(68),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_61: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(90),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(90),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_59: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(100),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(100),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_57: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(99),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(99),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_54: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(76),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(76),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_28: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(98),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(98),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_51: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(87),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(87),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_49: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(97),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(97),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_47: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(74),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(74),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_45: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(95),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(95),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_43: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(94),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(94),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_41: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(88),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(88),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_39: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(89),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(89),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_37: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(68),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(68),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_34: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(92),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(92),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_32: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(91),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(91),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_30: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(90),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(90),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_24: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(87),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(87),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_16: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_372__G1_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_372__G1\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_5: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(113),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(113),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_29: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_318__G1_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_318__G1\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_25: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_319__G1_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_319__G1\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_70: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_67: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_21: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_3_I_RETO\(0),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_3_I\(0),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_18: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0_RETO\(114),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(114),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_17: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1_RETO\(114),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(114),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_13: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0_RETO\(115),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(115),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_12: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1_RETO\(115),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(115),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_21: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3729_I_0\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_12: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(3),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT\(3),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_9: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(72),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(72),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_4: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(72),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(72),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_R_MK_BUSY_RET_8: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.BUSYMULXFF.UN2_TEMP_2_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.BUSYMULXFF.UN2_TEMP_2\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_R_MK_BUSY_RET_7: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3924_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3924\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_66: stratixii_lcell_ff port map (
regout => N_79941_RETO,
datain => N_79941,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RET_6: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_RETO\(9),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(9),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RET_5: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_RETO\(8),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(8),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RET_4: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.TEMP_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.TEMP\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RET_0: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.UN17_U_RDN_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.UN17_U_RDN\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RET_2: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.U_RDN_1_RETO\(1),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.U_RDN_1\(1),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RET: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_I_I_0_RETO\(0),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_I_I_0\(0),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_58: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RET_3: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RET_1: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_64: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(82),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_63: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(81),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_62: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_R_MK_BUSY_RET_1: stratixii_lcell_ff port map (
regout => RST_RETO,
datain => N_7,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_56: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2457_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2457\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_52: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_4_0_RETO\(4),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_4_0\(4),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_51: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2555_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2555\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_48: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_255_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_255\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_47: stratixii_lcell_ff port map (
regout => N_31723_1_RETO,
datain => N_31723_1,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_46: stratixii_lcell_ff port map (
regout => N_31763_1_RETO,
datain => N_31763_1,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_19: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5394\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5394_RETI\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_58_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(58),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(8),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(8),
clk => N_8,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_1: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10751_RETI\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G0_I_0\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G0_I_0_RETI\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_16_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(10),
clk => N_8,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(1),
clk => N_8,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_18: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349_I_0\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349_I_0_RETI\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_376_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(376),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_DIVMULTV\(0),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_14_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(14),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(14),
clk => N_8,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_45: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO(12),
datain => N_62,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_44: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO\(84),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M\(84),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_43: stratixii_lcell_ff port map (
regout => N_28952_RETO,
datain => N_28952,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_41: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO(8),
datain => N_58,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_40: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO\(6),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M\(6),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_39: stratixii_lcell_ff port map (
regout => N_28951_RETO,
datain => N_28951,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_37: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO(5),
datain => N_55,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_36: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO\(79),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M\(79),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_35: stratixii_lcell_ff port map (
regout => N_28950_RETO,
datain => N_28950,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_33: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO(10),
datain => N_60,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_32: stratixii_lcell_ff port map (
regout => N_28945_RETO,
datain => N_28945,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_31: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_29: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO(7),
datain => N_57,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_28: stratixii_lcell_ff port map (
regout => N_28947_RETO,
datain => N_28947,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_27: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO\(2),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M\(2),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_23: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO(11),
datain => N_61,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_17: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO(9),
datain => N_59,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_16: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_15: stratixii_lcell_ff port map (
regout => N_28946_RETO,
datain => N_28946,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_10: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_9: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(84),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_8: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_729_RETO\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_729\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_375_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(375),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(375),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_13_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(13),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(13),
clk => N_8,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_RETI\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_R_I_V: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.V\,
datain => N_48775,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_67_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(67),
datain => N_48774,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_R_I_RES_63_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(63),
datain => \GRLFPC2_0.COMB.V.I.RES_1\(63),
clk => N_8,
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_59_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(59),
datain => \GRLFPC2_0.FPO.EXP\(7),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(62),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_58_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(58),
datain => \GRLFPC2_0.FPO.EXP\(6),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(61),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_57_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(57),
datain => \GRLFPC2_0.FPO.EXP\(5),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(60),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_56_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(56),
datain => \GRLFPC2_0.FPO.EXP\(4),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(59),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_55_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(55),
datain => \GRLFPC2_0.FPO.EXP\(3),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(58),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_54_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(54),
datain => \GRLFPC2_0.FPO.EXP\(2),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(57),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_53_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(53),
datain => \GRLFPC2_0.FPO.EXP\(1),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(56),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_52_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(52),
datain => \GRLFPC2_0.FPO.EXP\(0),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(55),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_51_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(51),
datain => \GRLFPC2_0.FPO.FRAC\(54),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(54),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_50_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(50),
datain => \GRLFPC2_0.FPO.FRAC\(53),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(53),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_49_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(49),
datain => \GRLFPC2_0.FPO.FRAC\(52),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(52),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_48_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(48),
datain => \GRLFPC2_0.FPO.FRAC\(51),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(51),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_47_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(47),
datain => \GRLFPC2_0.FPO.FRAC\(50),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(50),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_46_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(46),
datain => \GRLFPC2_0.FPO.FRAC\(49),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(49),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_45_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(45),
datain => \GRLFPC2_0.FPO.FRAC\(48),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(48),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_44_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(44),
datain => \GRLFPC2_0.FPO.FRAC\(47),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(47),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_43_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(43),
datain => \GRLFPC2_0.FPO.FRAC\(46),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(46),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_42_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(42),
datain => \GRLFPC2_0.FPO.FRAC\(45),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(45),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_41_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(41),
datain => \GRLFPC2_0.FPO.FRAC\(44),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(44),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_40_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(40),
datain => \GRLFPC2_0.FPO.FRAC\(43),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(43),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_39_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(39),
datain => \GRLFPC2_0.FPO.FRAC\(42),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(42),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_38_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(38),
datain => \GRLFPC2_0.FPO.FRAC\(41),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(41),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_37_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(37),
datain => \GRLFPC2_0.FPO.FRAC\(40),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(40),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_36_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(36),
datain => \GRLFPC2_0.FPO.FRAC\(39),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(39),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_35_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(35),
datain => \GRLFPC2_0.FPO.FRAC\(38),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(38),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_34_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(34),
datain => \GRLFPC2_0.FPO.FRAC\(37),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(37),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_33_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(33),
datain => \GRLFPC2_0.FPO.FRAC\(36),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(36),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_32_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(32),
datain => \GRLFPC2_0.FPO.FRAC\(35),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(35),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_31_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(31),
datain => \GRLFPC2_0.FPO.FRAC\(34),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(34),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_30_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(30),
datain => \GRLFPC2_0.FPO.FRAC\(33),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(33),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_29_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(29),
datain => \GRLFPC2_0.FPO.FRAC\(32),
clk => N_8,
sload => \GRLFPC2_0.N_1470\,
adatasdata => \GRLFPC2_0.FPI.OP2\(32),
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_116_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(116),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2\,
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(118),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_117_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(117),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_175__G2\,
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(119),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_118_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(118),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_176__G2\,
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(120),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_119_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(119),
datain => \GRLFPC2_0.FPO.FRAC\(54),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(121),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_120_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(120),
datain => \GRLFPC2_0.FPO.FRAC\(53),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(122),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_121_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(121),
datain => \GRLFPC2_0.FPO.FRAC\(52),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(123),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_122_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(122),
datain => \GRLFPC2_0.FPO.FRAC\(51),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(124),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_123_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(123),
datain => \GRLFPC2_0.FPO.FRAC\(50),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(125),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_124_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(124),
datain => \GRLFPC2_0.FPO.FRAC\(49),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(126),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_125_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(125),
datain => \GRLFPC2_0.FPO.FRAC\(48),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(127),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_126_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(126),
datain => \GRLFPC2_0.FPO.FRAC\(47),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(128),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_127_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(127),
datain => \GRLFPC2_0.FPO.FRAC\(46),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(129),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_128_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(128),
datain => \GRLFPC2_0.FPO.FRAC\(45),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(130),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_129_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(129),
datain => \GRLFPC2_0.FPO.FRAC\(44),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(131),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_130_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(130),
datain => \GRLFPC2_0.FPO.FRAC\(43),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(132),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_131_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(131),
datain => \GRLFPC2_0.FPO.FRAC\(42),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(133),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_132_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(132),
datain => \GRLFPC2_0.FPO.FRAC\(41),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(134),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_133_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(133),
datain => \GRLFPC2_0.FPO.FRAC\(40),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(135),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_134_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(134),
datain => \GRLFPC2_0.FPO.FRAC\(39),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(136),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_135_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(135),
datain => \GRLFPC2_0.FPO.FRAC\(38),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(137),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_136_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(136),
datain => \GRLFPC2_0.FPO.FRAC\(37),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(138),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_137_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(137),
datain => \GRLFPC2_0.FPO.FRAC\(36),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(139),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_138_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(138),
datain => \GRLFPC2_0.FPO.FRAC\(35),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(140),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_139_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(139),
datain => \GRLFPC2_0.FPO.FRAC\(34),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(141),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_140_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(140),
datain => \GRLFPC2_0.FPO.FRAC\(33),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(142),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_141_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(141),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(141),
clk => N_8,
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_142_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(142),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(142),
clk => N_8,
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_143_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(143),
datain => \GRLFPC2_0.FPO.FRAC\(30),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(145),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_144_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(144),
datain => \GRLFPC2_0.FPO.FRAC\(29),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(146),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_145_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(145),
datain => \GRLFPC2_0.FPO.FRAC\(28),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(147),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_146_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(146),
datain => \GRLFPC2_0.FPO.FRAC\(27),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(148),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_147_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(147),
datain => \GRLFPC2_0.FPO.FRAC\(26),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(149),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_148_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(148),
datain => \GRLFPC2_0.FPO.FRAC\(25),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(150),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_149_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(149),
datain => \GRLFPC2_0.FPO.FRAC\(24),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(151),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_150_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(150),
datain => \GRLFPC2_0.FPO.FRAC\(23),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(152),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_151_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(151),
datain => \GRLFPC2_0.FPO.FRAC\(22),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(153),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_152_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(152),
datain => \GRLFPC2_0.FPO.FRAC\(21),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(154),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_153_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(153),
datain => \GRLFPC2_0.FPO.FRAC\(20),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(155),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_154_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(154),
datain => \GRLFPC2_0.FPO.FRAC\(19),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(156),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_155_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(155),
datain => \GRLFPC2_0.FPO.FRAC\(18),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(157),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_156_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(156),
datain => \GRLFPC2_0.FPO.FRAC\(17),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(158),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_157_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(157),
datain => \GRLFPC2_0.FPO.FRAC\(16),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(159),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_158_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(158),
datain => \GRLFPC2_0.FPO.FRAC\(15),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(160),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_159_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(159),
datain => \GRLFPC2_0.FPO.FRAC\(14),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(161),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_160_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(160),
datain => \GRLFPC2_0.FPO.FRAC\(13),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(162),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_161_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(161),
datain => \GRLFPC2_0.FPO.FRAC\(12),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(163),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_162_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(162),
datain => \GRLFPC2_0.FPO.FRAC\(11),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(164),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_163_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(163),
datain => \GRLFPC2_0.FPO.FRAC\(10),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(165),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_164_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(164),
datain => \GRLFPC2_0.FPO.FRAC\(9),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(166),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_165_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(165),
datain => \GRLFPC2_0.FPO.FRAC\(8),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(167),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_166_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(166),
datain => \GRLFPC2_0.FPO.FRAC\(7),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(168),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_167_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(167),
datain => \GRLFPC2_0.FPO.FRAC\(6),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(169),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_168_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(168),
datain => \GRLFPC2_0.FPO.FRAC\(5),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(170),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_169_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(169),
datain => \GRLFPC2_0.FPO.FRAC\(4),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(171),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_170_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(170),
datain => \GRLFPC2_0.FPO.FRAC\(3),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(172),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_171_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(171),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(2),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_14\(171),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_172_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(172),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(1),
clk => N_8,
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10381_I\,
adatasdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_14\(172),
ena => N_76337,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_247_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(247),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(247),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_248_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(248),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(248),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_249_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(249),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(249),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_250_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(250),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(250),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_251_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(251),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(251),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_252_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(252),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(252),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_253_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(253),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(253),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_254_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(254),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(254),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_255_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(255),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(255),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_256_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(256),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(256),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_257_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(257),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(257),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_77_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6_I\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_76_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(76),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7272\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_74_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(74),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7274\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_71_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(71),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.UN36_PCTRL_NEW_I\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_70_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(70),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(68),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_68_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(68),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3926\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_66_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(66),
datain => \GRLFPC2_0.FPI.START\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_65_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1780_I\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_64_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(64),
datain => \GRLFPC2_0.FPI.RST\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_63_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(63),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_62_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(62),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_61_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(61),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_60_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(60),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_59_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(59),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_58_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(58),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_57_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(57),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_56_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(56),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_55_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(55),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_54_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(54),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_53_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(53),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_52_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_51_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(51),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_50_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(50),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_49_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(49),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_48_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(48),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_48__I0_I_2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_47_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(47),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_47__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_46_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(46),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19\(45),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_45_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_44_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_44__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_43_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(43),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_43__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_42_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_41_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(41),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_41__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_40_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(40),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_40__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_39_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(39),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_39__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_38_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(38),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_16_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(16),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SCTRL_NEW\(0),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_15_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datain => N_81986,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_14_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(14),
datain => N_59162,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_13_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(13),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7248\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_12_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(12),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_I_I_0\(0),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_11_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datain => N_81985,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_10_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_9_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(9),
datain => N_35958,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.TEMP\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_8_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(8),
datain => N_35959,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.TEMP\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_6_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(6),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4459\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_5_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(5),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_2_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(2),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7259\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_1_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(1),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7260\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(0),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW_6\(0),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_36_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_35_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(35),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_35__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_34_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_33_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_32_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_31_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__I0_I_0\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_30_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_30__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_29_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_28_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_27_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_26_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_25_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_24_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(24),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_24__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_23_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(23),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_23__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_22_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(22),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_22__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_21_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(21),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_21__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_20_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(20),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_20__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_19_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(19),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_18_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(18),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(5),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(2),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_2__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(1),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_1__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_377_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(377),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(0),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_373_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(373),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_3_I\(0),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_372_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(372),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_372__G1\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_371_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(371),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(112),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_370_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(370),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(111),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_369_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(369),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(110),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_368_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(368),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(109),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_367_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(367),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(108),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_366_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(366),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(107),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_365_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(365),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(106),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_364_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(364),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(105),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_363_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(363),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(104),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_362_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(362),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(103),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_361_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(361),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(102),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_360_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(360),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(101),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_359_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(359),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(100),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_358_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(358),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(99),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_357_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(357),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(98),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_356_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(356),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(97),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_355_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(355),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(96),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_354_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(354),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(95),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_353_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(353),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(94),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_352_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(352),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(93),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_351_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(351),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(92),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_350_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(350),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(91),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_349_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(349),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(90),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_348_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(348),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(89),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_347_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(347),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(88),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_346_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(346),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(87),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_345_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(345),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(86),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_344_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(344),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(85),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_343_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(343),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(84),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_342_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(342),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(83),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_341_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(341),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(82),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_340_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(340),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(81),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_339_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(339),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(80),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_338_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(338),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(79),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_337_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(337),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(78),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_336_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(336),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(77),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_335_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(335),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(76),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_334_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(334),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(75),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_333_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(333),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(74),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_332_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(332),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(73),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_331_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(331),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(72),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_330_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(330),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(71),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_329_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(329),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(70),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_328_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(328),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(69),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_327_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(327),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(68),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_326_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(326),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(67),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_325_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(325),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(66),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_324_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(324),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(65),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_323_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(323),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(64),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_322_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(322),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(63),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_321_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(321),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(62),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_320_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(320),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(61),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_319_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(319),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_319__G1\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_318_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(318),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_318__G1\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_317_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(317),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_317__G1\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_316_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(316),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_316__G1\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_315_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(315),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_314_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(314),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(55),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_313_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(313),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(54),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_312_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(312),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(53),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_311_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(311),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(52),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_310_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(310),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(51),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_309_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(309),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(50),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_308_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(308),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(49),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_307_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(307),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(48),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_306_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(306),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(47),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_305_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(305),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(46),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_304_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(304),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(45),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_303_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(303),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(44),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_302_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(302),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(43),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_301_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(301),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(42),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_300_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(300),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(41),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_299_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(299),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(40),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_298_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(298),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(39),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_297_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(297),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(38),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_296_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(296),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(37),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_295_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(295),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(36),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_294_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(294),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(35),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_293_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(293),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(34),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_292_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(292),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(33),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_291_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(291),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(32),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_290_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(290),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(31),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_289_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(289),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(30),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_288_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(288),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(29),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_287_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(287),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(28),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_286_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(286),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(27),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_285_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(285),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(26),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_284_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(284),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(25),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_283_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(283),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(24),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_282_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(282),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(23),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_281_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(281),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(22),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_280_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(280),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(21),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_279_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(279),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(20),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_278_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(278),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(19),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_277_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(277),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(18),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_276_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(276),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(17),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_275_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(275),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(16),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_274_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(274),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(15),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_273_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(273),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(14),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_272_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(272),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(13),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_271_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(271),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(12),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_270_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(270),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(11),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_269_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(269),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(10),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_268_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(268),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(9),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_267_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(267),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(8),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_266_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(266),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(7),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_265_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(265),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(6),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_264_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(264),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(5),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_263_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(263),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(4),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_262_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(262),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(3),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_261_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(261),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(2),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_260_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(260),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(1),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_259_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(259),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(0),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_258_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(258),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_258__N_5_I\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_246_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(246),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_245_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(245),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(245),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_244_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244),
datain => N_36366,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_243_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(243),
datain => N_36367,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_242_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242),
datain => N_36368,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_241_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(241),
datain => N_36369,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_240_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(240),
datain => N_36370,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_239_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(239),
datain => N_36371,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_238_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(238),
datain => N_36372,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_237_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(237),
datain => N_36373,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_236_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236),
datain => N_36149,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_235_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235),
datain => N_36176,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_234_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234),
datain => N_36203,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_233_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233),
datain => N_36374,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_232_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(232),
datain => N_36375,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_230_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(230),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(1),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_229_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(229),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(2),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_228_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(228),
datain => \GRLFPC2_0.FPO.FRAC\(3),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_227_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(227),
datain => \GRLFPC2_0.FPO.FRAC\(4),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_226_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(226),
datain => \GRLFPC2_0.FPO.FRAC\(5),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_225_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(225),
datain => \GRLFPC2_0.FPO.FRAC\(6),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_224_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(224),
datain => \GRLFPC2_0.FPO.FRAC\(7),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_223_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(223),
datain => \GRLFPC2_0.FPO.FRAC\(8),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_222_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(222),
datain => \GRLFPC2_0.FPO.FRAC\(9),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_221_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(221),
datain => \GRLFPC2_0.FPO.FRAC\(10),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_220_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(220),
datain => \GRLFPC2_0.FPO.FRAC\(11),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_219_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(219),
datain => \GRLFPC2_0.FPO.FRAC\(12),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_218_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(218),
datain => \GRLFPC2_0.FPO.FRAC\(13),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_217_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(217),
datain => \GRLFPC2_0.FPO.FRAC\(14),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_216_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(216),
datain => \GRLFPC2_0.FPO.FRAC\(15),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_215_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(215),
datain => \GRLFPC2_0.FPO.FRAC\(16),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_214_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(214),
datain => \GRLFPC2_0.FPO.FRAC\(17),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_213_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(213),
datain => \GRLFPC2_0.FPO.FRAC\(18),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_212_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(212),
datain => \GRLFPC2_0.FPO.FRAC\(19),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_211_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(211),
datain => \GRLFPC2_0.FPO.FRAC\(20),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_210_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(210),
datain => \GRLFPC2_0.FPO.FRAC\(21),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_209_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(209),
datain => \GRLFPC2_0.FPO.FRAC\(22),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_208_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(208),
datain => \GRLFPC2_0.FPO.FRAC\(23),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_207_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(207),
datain => \GRLFPC2_0.FPO.FRAC\(24),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_206_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(206),
datain => \GRLFPC2_0.FPO.FRAC\(25),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_205_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(205),
datain => \GRLFPC2_0.FPO.FRAC\(26),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_204_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(204),
datain => \GRLFPC2_0.FPO.FRAC\(27),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_203_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(203),
datain => \GRLFPC2_0.FPO.FRAC\(28),
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_202_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(202),
datain => N_26536,
clk => N_8,
sload => N_26534_I,
adatasdata => N_26535,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
N_26534_I <= not N_26534;
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_201_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(201),
datain => N_26538,
clk => N_8,
sload => N_26534_I,
adatasdata => N_26537,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_200_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(200),
datain => N_26540,
clk => N_8,
sload => N_26534_I,
adatasdata => N_26539,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_199_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(199),
datain => N_26542,
clk => N_8,
sload => N_26534_I,
adatasdata => N_26541,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_198_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(198),
datain => N_26544,
clk => N_8,
sload => N_26534_I,
adatasdata => N_26543,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_197_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(197),
datain => N_26546,
clk => N_8,
sload => N_26534_I,
adatasdata => N_26545,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_196_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(196),
datain => N_26548,
clk => N_8,
sload => N_26534_I,
adatasdata => N_26547,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_195_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(195),
datain => N_26550,
clk => N_8,
sload => N_26534_I,
adatasdata => N_26549,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_194_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(194),
datain => N_26552,
clk => N_8,
sload => N_26534_I,
adatasdata => N_26551,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_193_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(193),
datain => N_26554,
clk => N_8,
sload => N_26534_I,
adatasdata => N_26553,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_192_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(192),
datain => N_26556,
clk => N_8,
sload => N_26534_I,
adatasdata => N_26555,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_191_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(191),
datain => N_26558,
clk => N_8,
sload => N_26534_I,
adatasdata => N_26557,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_190_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(190),
datain => N_26560,
clk => N_8,
sload => N_26534_I,
adatasdata => N_26559,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_189_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(189),
datain => N_26562,
clk => N_8,
sload => N_26534_I,
adatasdata => N_26561,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_188_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(188),
datain => N_26564,
clk => N_8,
sload => N_26534_I,
adatasdata => N_26563,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_187_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(187),
datain => N_26566,
clk => N_8,
sload => N_26534_I,
adatasdata => N_26565,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_186_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(186),
datain => N_26568,
clk => N_8,
sload => N_26534_I,
adatasdata => N_26567,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_185_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(185),
datain => N_26570,
clk => N_8,
sload => N_26534_I,
adatasdata => N_26569,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_184_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(184),
datain => N_26572,
clk => N_8,
sload => N_26534_I,
adatasdata => N_26571,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_183_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(183),
datain => N_26574,
clk => N_8,
sload => N_26534_I,
adatasdata => N_26573,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_182_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(182),
datain => N_26576,
clk => N_8,
sload => N_26534_I,
adatasdata => N_26575,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_181_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(181),
datain => N_26578,
clk => N_8,
sload => N_26534_I,
adatasdata => N_26577,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_180_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(180),
datain => N_26580,
clk => N_8,
sload => N_26534_I,
adatasdata => N_26579,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_179_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(179),
datain => N_26582,
clk => N_8,
sload => N_26534_I,
adatasdata => N_26581,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_178_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(178),
datain => N_26584,
clk => N_8,
sload => N_26534_I,
adatasdata => N_26583,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_177_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(177),
datain => N_26586,
clk => N_8,
sload => N_26534_I,
adatasdata => N_26585,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_176_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(176),
datain => N_26588,
clk => N_8,
sload => N_26534_I,
adatasdata => N_26587,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_175_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(175),
datain => N_26590,
clk => N_8,
sload => N_26534_I,
adatasdata => N_26589,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_174_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(174),
datain => N_26592,
clk => N_8,
sload => N_26534_I,
adatasdata => N_26591,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_173_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(173),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(173),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_R_MK_HOLDN2: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.MK.HOLDN2\,
datain => \GRLFPC2_0.R.MK.HOLDN1\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_R_MK_RST2: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.MK.RST2\,
datain => \GRLFPC2_0.R.MK.RST\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_R_MK_RST_RET: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.COMB.ANNULFPU_1_O\,
datain => \GRLFPC2_0.COMB.ANNULFPU_1\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_R_MK_RST_RET_6: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.MK.HOLDN2_O\,
datain => \GRLFPC2_0.R.MK.HOLDN2\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_R_MK_RST_RET_2: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.MK.RST2_O\,
datain => \GRLFPC2_0.R.MK.RST2\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_R_MK_LDOP_RET: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.HOLDN_O\,
datain => N_9,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_R_MK_LDOP_RET_3: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.COMB.LOCKGEN.LOCKI_O_3\,
datain => \GRLFPC2_0.COMB.LOCKGEN.LOCKI_I_I\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_R_MK_LDOP_RET_6: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O_3\(0),
datain => N_10,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_R_M_AFQ_RET_1: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.N_1829_O\,
datain => \GRLFPC2_0.N_1683\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_E_AFQ_RET_1: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.N_1830_O\,
datain => \GRLFPC2_0.N_1237\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_M_AFQ_RET: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.E.AFQ_O\,
datain => \GRLFPC2_0.R.M.AFQ_RET_0_0_G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_M_AFSR_RET: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.E.AFSR_O\,
datain => \GRLFPC2_0.R.M.AFSR_RET_0_0_G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_A_RS2D: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.A.RS2D\,
datain => \GRLFPC2_0.COMB.RS2D_1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_A_RS1D: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.A.RS1D\,
datain => \GRLFPC2_0.COMB.RS1D_1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_M_SEQERR: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.N_554\,
datain => \GRLFPC2_0.N_553\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_A_SEQERR_RET_3: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.N_1837_O\,
datain => \GRLFPC2_0.N_835\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_A_AFQ_RET_5: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(0),
datain => N_10,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_E_AFQ_RET: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.A.AFQ_O\,
datain => \GRLFPC2_0.R.A.AFQ\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_A_ST_RET: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.COMB.FPDECODE.ST_O\,
datain => \GRLFPC2_0.COMB.FPDECODE.ST\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_E_SEQERR: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.N_553\,
datain => \GRLFPC2_0.R.E.SEQERR_0_0_G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_E_AFSR_RET: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.A.AFSR_O\,
datain => \GRLFPC2_0.R.A.AFSR\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_I_PC_RET_60: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datain => \GRLFPC2_0.V.I.EXEC_0_SQMUXA\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_A_AFQ_RET_2: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.COMB.LOCKGEN.LOCKI_O\,
datain => \GRLFPC2_0.COMB.LOCKGEN.LOCKI_I_I\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_X_RDD: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.X.RDD\,
datain => \GRLFPC2_0.N_559\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_M_RDD: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.N_559\,
datain => \GRLFPC2_0.N_558\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_E_RDD: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.N_558\,
datain => \GRLFPC2_0.N_557\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_A_RDD: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.N_557\,
datain => \GRLFPC2_0.R.A.RDD_0_0_G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_X_SEQERR: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.X.SEQERR\,
datain => \GRLFPC2_0.N_554\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_A_LD: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.A.LD\,
datain => \GRLFPC2_0.R.A.LD_0_0_G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_A_FPOP: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.A.FPOP\,
datain => \GRLFPC2_0.N_1000\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
RST_I <= not N_7;
GRLFPC2_0_R_I_EXEC: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.EXEC\,
datain => \GRLFPC2_0.COMB.V.I.EXEC_1_3\,
clk => N_8,
sclr => RST_I,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_FSR_FTT_2_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.FSR.FTT\(2),
datain => \GRLFPC2_0.N_50_1\,
clk => N_8,
sclr => RST_I,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_FSR_FTT_0_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.FSR.FTT\(0),
datain => \GRLFPC2_0.R.FSR.FTT_0_0_0__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_FSR_NONSTD: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.FSR.NONSTD\,
datain => \GRLFPC2_0.R.FSR.NONSTD_0_0_G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_I_RDD: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RDD\,
datain => \GRLFPC2_0.R.I.RDD_0_0_G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_X_LD: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.X.LD\,
datain => \GRLFPC2_0.R.X.LD_0_0_G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_X_FPOP: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.X.FPOP\,
datain => \GRLFPC2_0.R.X.FPOP_0_0_G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_X_AFSR: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.X.AFSR\,
datain => \GRLFPC2_0.R.X.AFSR_0_0_G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_X_AFQ: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.X.AFQ\,
datain => \GRLFPC2_0.R.X.AFQ_0_0_G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_M_LD: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.M.LD\,
datain => \GRLFPC2_0.R.M.LD_0_0_G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_M_FPOP: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.M.FPOP\,
datain => \GRLFPC2_0.R.M.FPOP_0_0_G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_E_LD: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.E.LD\,
datain => \GRLFPC2_0.R.E.LD_0_0_G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_E_FPOP: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.E.FPOP\,
datain => \GRLFPC2_0.COMB.V.E.FPOP_1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_R_MK_HOLDN1: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.MK.HOLDN1\,
datain => \GRLFPC2_0.N_2101\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_R_MK_BUSY2_RET: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.COMB.ANNULFPU_1_O_0\,
datain => \GRLFPC2_0.COMB.ANNULFPU_1\,
clk => N_8,
sclr => RST_I,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_R_MK_BUSY_RET_3: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.MK.HOLDN2_O_0\,
datain => \GRLFPC2_0.R.MK.HOLDN2\,
clk => N_8,
sclr => RST_I,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_R_MK_BUSY_RET_2: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.MK.HOLDN1_O_0\,
datain => \GRLFPC2_0.R.MK.HOLDN1\,
clk => N_8,
sclr => RST_I,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_R_MK_BUSY2_RET_1: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.MK.BUSY_O\,
datain => \GRLFPC2_0.N_2111\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_R_MK_BUSY_RET_5: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.MK.RST2_O_0\,
datain => \GRLFPC2_0.R.MK.RST2\,
clk => N_8,
sclr => RST_I,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_R_MK_BUSY_RET_4: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.MK.RST_O_0\,
datain => \GRLFPC2_0.N_2115\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_R_I_INST_0_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(0),
datain => N_326,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_1_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(1),
datain => N_327,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_2_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(2),
datain => N_328,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_3_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(3),
datain => N_329,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_4_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(4),
datain => N_330,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_5_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(5),
datain => N_331,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_6_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(6),
datain => N_332,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_7_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(7),
datain => N_333,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_8_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(8),
datain => N_334,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_9_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(9),
datain => N_335,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_10_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(10),
datain => N_336,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_11_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(11),
datain => N_337,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_12_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(12),
datain => N_338,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_13_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(13),
datain => N_339,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_14_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(14),
datain => N_340,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_15_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(15),
datain => N_341,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_16_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(16),
datain => N_342,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_17_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(17),
datain => N_343,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_18_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(18),
datain => N_344,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_19_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(19),
datain => N_345,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_20_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(20),
datain => N_346,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_21_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(21),
datain => N_347,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_22_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(22),
datain => N_348,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_23_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(23),
datain => N_349,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_24_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(24),
datain => N_350,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_25_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(25),
datain => N_351,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_26_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(26),
datain => N_352,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_27_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(27),
datain => N_353,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_28_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(28),
datain => N_354,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_29_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(29),
datain => N_355,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_30_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(30),
datain => N_356,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_INST_31_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.INST\(31),
datain => N_357,
clk => N_8,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_0_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(0),
datain => \GRLFPC2_0.R.E.STDATA_1_0_0__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_1_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(1),
datain => \GRLFPC2_0.R.E.STDATA_1_0_1__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_2_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(2),
datain => \GRLFPC2_0.R.E.STDATA_1_0_2__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_3_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(3),
datain => \GRLFPC2_0.R.E.STDATA_1_0_3__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_4_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(4),
datain => \GRLFPC2_0.R.E.STDATA_1_0_4__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_5_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(5),
datain => \GRLFPC2_0.R.E.STDATA_1_0_5__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_6_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(6),
datain => \GRLFPC2_0.R.E.STDATA_1_0_6__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_7_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(7),
datain => \GRLFPC2_0.R.E.STDATA_1_0_7__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_8_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(8),
datain => \GRLFPC2_0.R.E.STDATA_1_0_8__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_9_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(9),
datain => \GRLFPC2_0.R.E.STDATA_1_0_9__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_10_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(10),
datain => \GRLFPC2_0.R.E.STDATA_1_0_10__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_11_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(11),
datain => \GRLFPC2_0.R.E.STDATA_1_0_11__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_12_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(12),
datain => \GRLFPC2_0.R.E.STDATA_1_0_12__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_13_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(13),
datain => \GRLFPC2_0.R.E.STDATA_1_0_13__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_14_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(14),
datain => \GRLFPC2_0.R.E.STDATA_1_0_14__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_15_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(15),
datain => \GRLFPC2_0.R.E.STDATA_1_0_15__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_16_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(16),
datain => \GRLFPC2_0.R.E.STDATA_1_0_16__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_17_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(17),
datain => \GRLFPC2_0.R.E.STDATA_1_0_17__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_18_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(18),
datain => \GRLFPC2_0.R.E.STDATA_1_0_18__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_19_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(19),
datain => \GRLFPC2_0.R.E.STDATA_1_0_19__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_20_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(20),
datain => \GRLFPC2_0.R.E.STDATA_1_0_20__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_21_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(21),
datain => \GRLFPC2_0.R.E.STDATA_1_0_21__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_22_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(22),
datain => \GRLFPC2_0.R.E.STDATA_1_0_22__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_23_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(23),
datain => \GRLFPC2_0.R.E.STDATA_1_0_23__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_24_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(24),
datain => \GRLFPC2_0.R.E.STDATA_1_0_24__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_25_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(25),
datain => \GRLFPC2_0.R.E.STDATA_1_0_25__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_26_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(26),
datain => \GRLFPC2_0.R.E.STDATA_1_0_26__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_27_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(27),
datain => \GRLFPC2_0.R.E.STDATA_1_0_27__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_28_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(28),
datain => \GRLFPC2_0.R.E.STDATA_1_0_28__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_29_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(29),
datain => \GRLFPC2_0.R.E.STDATA_1_0_29__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_30_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(30),
datain => \GRLFPC2_0.R.E.STDATA_1_0_30__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_E_STDATA_31_\: stratixii_lcell_ff port map (
regout => CPO_DATAZ(31),
datain => \GRLFPC2_0.R.E.STDATA_1_0_31__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_FSR_RD_0_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.FSR.RD\(0),
datain => \GRLFPC2_0.R.FSR.RD_0_0_0__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_FSR_RD_1_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.FSR.RD\(1),
datain => \GRLFPC2_0.R.FSR.RD_0_0_1__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_FSR_TEM_0_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.FSR.TEM\(0),
datain => \GRLFPC2_0.R.FSR.TEM_1_0_0__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_FSR_TEM_1_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.FSR.TEM\(1),
datain => \GRLFPC2_0.R.FSR.TEM_1_0_1__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_FSR_TEM_2_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.FSR.TEM\(2),
datain => \GRLFPC2_0.R.FSR.TEM_1_0_2__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_FSR_TEM_3_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.FSR.TEM\(3),
datain => \GRLFPC2_0.R.FSR.TEM_1_0_3__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_FSR_TEM_4_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.FSR.TEM\(4),
datain => \GRLFPC2_0.R.FSR.TEM_1_0_4__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_STATE_0_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.STATE\(0),
datain => \GRLFPC2_0.R.STATE_0_0_0__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_STATE_1_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.STATE\(1),
datain => \GRLFPC2_0.R.STATE_0_0_1__I0_I_1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_A_RF1REN_2_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.A.RF1REN\(2),
datain => N_36379,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_A_RF1REN_1_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.A.RF1REN\(1),
datain => N_36380,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_A_RF2REN_2_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.A.RF2REN\(2),
datain => N_36381,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_A_RF2REN_1_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.A.RF2REN\(1),
datain => N_36382,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_FSR_FCC_0_\: stratixii_lcell_ff port map (
regout => CPO_CCZ(0),
datain => \GRLFPC2_0.R.FSR.FCC_0_0_0__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_FSR_FCC_1_\: stratixii_lcell_ff port map (
regout => CPO_CCZ(1),
datain => \GRLFPC2_0.R.FSR.FCC_0_0_1__G1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_FSR_AEXC_0_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.FSR.AEXC\(0),
datain => \GRLFPC2_0.R.FSR.AEXC_1_0_0__I0_I_0\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_FSR_AEXC_1_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.FSR.AEXC\(1),
datain => \GRLFPC2_0.R.FSR.AEXC_1_0_1__I0_I_1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_FSR_AEXC_2_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.FSR.AEXC\(2),
datain => \GRLFPC2_0.R.FSR.AEXC_1_0_2__I0_I_0\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_FSR_AEXC_3_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.FSR.AEXC\(3),
datain => \GRLFPC2_0.R.FSR.AEXC_1_0_3__I0_I_1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_FSR_AEXC_4_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.FSR.AEXC\(4),
datain => \GRLFPC2_0.R.FSR.AEXC_1_0_4__I0_I_0\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_FSR_CEXC_0_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.FSR.CEXC\(0),
datain => \GRLFPC2_0.R.FSR.CEXC_1_0_0__I0_I_1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_FSR_CEXC_1_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.FSR.CEXC\(1),
datain => \GRLFPC2_0.R.FSR.CEXC_1_0_1__I0_I_0\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_FSR_CEXC_2_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.FSR.CEXC\(2),
datain => \GRLFPC2_0.R.FSR.CEXC_1_0_2__I0_I_1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_FSR_CEXC_3_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.FSR.CEXC\(3),
datain => \GRLFPC2_0.R.FSR.CEXC_1_0_3__I0_I_0\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_FSR_CEXC_4_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.FSR.CEXC\(4),
datain => \GRLFPC2_0.R.FSR.CEXC_1_0_4__I0_I_1\,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_A_MOV_RET_0_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(69),
datain => N_80,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_A_MOV_RET_2_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(44),
datain => N_55,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_A_MOV_RET_3_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(45),
datain => N_56,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_A_MOV_RET_4_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(46),
datain => N_57,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_A_MOV_RET_5_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(47),
datain => N_58,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_A_MOV_RET_6_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(48),
datain => N_59,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_A_MOV_RET_7_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(49),
datain => N_60,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_A_MOV_RET_8_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(50),
datain => N_61,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_A_MOV_RET_9_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(51),
datain => N_62,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_A_MOV_RET_10_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(52),
datain => N_63,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_A_MOV_RET_12_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(59),
datain => N_70,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_A_MOV_RET_15_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(62),
datain => N_73,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_A_SEQERR_RET_4_0_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.STATE_O\(0),
datain => \GRLFPC2_0.R.STATE\(0),
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_A_SEQERR_RET_4_1_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.STATE_O\(1),
datain => \GRLFPC2_0.R.STATE\(1),
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_A_AFQ_RET_0_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(73),
datain => N_84,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_A_AFQ_RET_1_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(74),
datain => N_85,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_A_AFQ_RET_2_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(58),
datain => N_69,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_A_AFQ_RET_4_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(60),
datain => N_71,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_A_AFQ_RET_5_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(61),
datain => N_72,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_A_AFQ_RET_7_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(63),
datain => N_74,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_A_AFQ_RET_9_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(70),
datain => N_81,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_CC_0_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.CC\(0),
datain => \GRLFPC2_0.R.I.CC_0_0_0__G2\,
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_CC_1_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.CC\(1),
datain => \GRLFPC2_0.R.I.CC_0_0_1__G2\,
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_0_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(2),
datain => \GRLFPC2_0.FPCI_O\(285),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_1_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(3),
datain => \GRLFPC2_0.FPCI_O\(286),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_2_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(4),
datain => \GRLFPC2_0.FPCI_O\(287),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_3_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(5),
datain => \GRLFPC2_0.FPCI_O\(288),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_4_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(6),
datain => \GRLFPC2_0.FPCI_O\(289),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_5_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(7),
datain => \GRLFPC2_0.FPCI_O\(290),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_6_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(8),
datain => \GRLFPC2_0.FPCI_O\(291),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_7_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(9),
datain => \GRLFPC2_0.FPCI_O\(292),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_8_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(10),
datain => \GRLFPC2_0.FPCI_O\(293),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_9_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(11),
datain => \GRLFPC2_0.FPCI_O\(294),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_10_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(12),
datain => \GRLFPC2_0.FPCI_O\(295),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_11_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(13),
datain => \GRLFPC2_0.FPCI_O\(296),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_12_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(14),
datain => \GRLFPC2_0.FPCI_O\(297),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_13_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(15),
datain => \GRLFPC2_0.FPCI_O\(298),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_14_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(16),
datain => \GRLFPC2_0.FPCI_O\(299),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_15_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(17),
datain => \GRLFPC2_0.FPCI_O\(300),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_16_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(18),
datain => \GRLFPC2_0.FPCI_O\(301),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_17_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(19),
datain => \GRLFPC2_0.FPCI_O\(302),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_18_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(20),
datain => \GRLFPC2_0.FPCI_O\(303),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_19_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(21),
datain => \GRLFPC2_0.FPCI_O\(304),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_20_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(22),
datain => \GRLFPC2_0.FPCI_O\(305),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_21_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(23),
datain => \GRLFPC2_0.FPCI_O\(306),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_22_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(24),
datain => \GRLFPC2_0.FPCI_O\(307),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_23_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(25),
datain => \GRLFPC2_0.FPCI_O\(308),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_24_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(26),
datain => \GRLFPC2_0.FPCI_O\(309),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_25_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(27),
datain => \GRLFPC2_0.FPCI_O\(310),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_26_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(28),
datain => \GRLFPC2_0.FPCI_O\(311),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_27_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(29),
datain => \GRLFPC2_0.FPCI_O\(312),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_28_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(30),
datain => \GRLFPC2_0.FPCI_O\(313),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_29_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.PC_O\(31),
datain => \GRLFPC2_0.FPCI_O\(314),
clk => N_8,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_0_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(285),
datain => N_296,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_1_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(286),
datain => N_297,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_2_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(287),
datain => N_298,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_3_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(288),
datain => N_299,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_4_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(289),
datain => N_300,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_5_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(290),
datain => N_301,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_6_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(291),
datain => N_302,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_7_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(292),
datain => N_303,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_8_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(293),
datain => N_304,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_9_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(294),
datain => N_305,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_10_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(295),
datain => N_306,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_11_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(296),
datain => N_307,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_12_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(297),
datain => N_308,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_13_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(298),
datain => N_309,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_14_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(299),
datain => N_310,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_15_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(300),
datain => N_311,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_16_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(301),
datain => N_312,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_17_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(302),
datain => N_313,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_18_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(303),
datain => N_314,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_19_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(304),
datain => N_315,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_20_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(305),
datain => N_316,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_21_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(306),
datain => N_317,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_22_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(307),
datain => N_318,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_23_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(308),
datain => N_319,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_24_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(309),
datain => N_320,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_25_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(310),
datain => N_321,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_26_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(311),
datain => N_322,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_27_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(312),
datain => N_323,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_28_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(313),
datain => N_324,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_PC_RET_30_29_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O\(314),
datain => N_325,
clk => N_8,
ena => N_9,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_EXC_0_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.EXC\(0),
datain => \GRLFPC2_0.R.I.EXC_MB\(0),
clk => N_8,
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_EXC_1_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.EXC\(1),
datain => \GRLFPC2_0.R.I.EXC_2_0_1__G2\,
clk => N_8,
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_EXC_2_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.EXC\(2),
datain => \GRLFPC2_0.R.I.EXC_2_0_2__G2\,
clk => N_8,
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_EXC_3_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.EXC\(3),
datain => \GRLFPC2_0.R.I.EXC_2_0_3__G2\,
clk => N_8,
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_EXC_4_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.EXC\(4),
datain => \GRLFPC2_0.R.I.EXC_2_0_4__G2\,
clk => N_8,
ena => \GRLFPC2_0.R.I.EXC_2_0_4__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_MK_LDOP_RET_4_0_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.STATE_O_3\(0),
datain => \GRLFPC2_0.R.STATE\(0),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_R_MK_LDOP_RET_4_1_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.STATE_O_3\(1),
datain => \GRLFPC2_0.R.STATE\(1),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_R_MK_LDOP_RET_1_0_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O_3\(73),
datain => N_84,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_R_MK_LDOP_RET_1_1_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O_3\(74),
datain => N_85,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_R_MK_LDOP_RET_1_2_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O_0\(63),
datain => N_74,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_R_MK_LDOP_RET_1_3_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O_0\(62),
datain => N_73,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_R_MK_LDOP_RET_1_4_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O_0\(61),
datain => N_72,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_R_MK_LDOP_RET_1_5_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O_0\(60),
datain => N_71,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_R_MK_LDOP_RET_1_6_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O_0\(59),
datain => N_70,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_R_MK_LDOP_RET_1_7_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O_0\(69),
datain => N_80,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_R_MK_LDOP_RET_1_8_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPCI_O_0\(70),
datain => N_81,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_R_A_RS1_0_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.A.RS1\(0),
datain => \GRLFPC2_0.COMB.RS1_1\(0),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_R_A_RS1_1_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.A.RS1\(1),
datain => \GRLFPC2_0.COMB.RS1_1\(1),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_R_A_RS1_2_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.A.RS1\(2),
datain => \GRLFPC2_0.COMB.RS1_1\(2),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_R_A_RS1_3_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.A.RS1\(3),
datain => \GRLFPC2_0.COMB.RS1_1\(3),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_R_A_RS1_4_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.A.RS1\(4),
datain => \GRLFPC2_0.COMB.RS1_1\(4),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_R_I_RES_0_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(0),
datain => \GRLFPC2_0.FPO.FRAC\(3),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_1_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(1),
datain => \GRLFPC2_0.FPO.FRAC\(4),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_2_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(2),
datain => \GRLFPC2_0.FPO.FRAC\(5),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_3_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(3),
datain => \GRLFPC2_0.FPO.FRAC\(6),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_4_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(4),
datain => \GRLFPC2_0.FPO.FRAC\(7),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_5_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(5),
datain => \GRLFPC2_0.FPO.FRAC\(8),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_6_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(6),
datain => \GRLFPC2_0.FPO.FRAC\(9),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_7_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(7),
datain => \GRLFPC2_0.FPO.FRAC\(10),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_8_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(8),
datain => \GRLFPC2_0.FPO.FRAC\(11),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_9_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(9),
datain => \GRLFPC2_0.FPO.FRAC\(12),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_10_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(10),
datain => \GRLFPC2_0.FPO.FRAC\(13),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_11_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(11),
datain => \GRLFPC2_0.FPO.FRAC\(14),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_12_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(12),
datain => \GRLFPC2_0.FPO.FRAC\(15),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_13_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(13),
datain => \GRLFPC2_0.FPO.FRAC\(16),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_14_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(14),
datain => \GRLFPC2_0.FPO.FRAC\(17),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_15_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(15),
datain => \GRLFPC2_0.FPO.FRAC\(18),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_16_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(16),
datain => \GRLFPC2_0.FPO.FRAC\(19),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_17_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(17),
datain => \GRLFPC2_0.FPO.FRAC\(20),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_18_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(18),
datain => \GRLFPC2_0.FPO.FRAC\(21),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_19_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(19),
datain => \GRLFPC2_0.FPO.FRAC\(22),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_20_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(20),
datain => \GRLFPC2_0.FPO.FRAC\(23),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_21_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(21),
datain => \GRLFPC2_0.FPO.FRAC\(24),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_22_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(22),
datain => \GRLFPC2_0.FPO.FRAC\(25),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_23_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(23),
datain => \GRLFPC2_0.FPO.FRAC\(26),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_24_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(24),
datain => \GRLFPC2_0.FPO.FRAC\(27),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_25_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(25),
datain => \GRLFPC2_0.FPO.FRAC\(28),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_26_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(26),
datain => \GRLFPC2_0.FPO.FRAC\(29),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_27_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(27),
datain => \GRLFPC2_0.FPO.FRAC\(30),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_28_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(28),
datain => \GRLFPC2_0.FPO.FRAC\(31),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_60_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(60),
datain => \GRLFPC2_0.FPO.EXP\(8),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_61_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(61),
datain => \GRLFPC2_0.FPO.EXP\(9),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_I_RES_62_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.I.RES\(62),
datain => \GRLFPC2_0.FPO.EXP\(10),
clk => N_8,
ena => \GRLFPC2_0.N_1255\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_R_A_RS2_0_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.A.RS2\(0),
datain => \GRLFPC2_0.COMB.RS2_1\(0),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_R_A_RS2_1_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.A.RS2\(1),
datain => \GRLFPC2_0.COMB.RS2_1\(1),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_R_A_RS2_2_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.A.RS2\(2),
datain => \GRLFPC2_0.COMB.RS2_1\(2),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_R_A_RS2_3_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.A.RS2\(3),
datain => \GRLFPC2_0.COMB.RS2_1\(3),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_R_A_RS2_4_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.R.A.RS2\(4),
datain => \GRLFPC2_0.COMB.RS2_1\(4),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_17_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_1\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_RNO_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_8\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_9\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1937\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2581\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2063\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1941\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_17_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_4\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_RNO_17_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_8\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_9\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1937\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2581\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2063\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1941\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_10_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_0\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIHTQC5_0_20_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"f0f05041f0f05050")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(20),
datae => \GRLFPC2_0.FPI.LDOP_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6_I\,
datac => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_42_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(42),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2_0\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_RNO_42_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcccf000ffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2_0\,
dataf => N_79943,
datae => N_32619_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2776\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2490\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3_0\(41));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_130: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_RETI_0\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNI02EQ71_16_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"faaaf000feeefccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_RETI_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(375),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_16_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI_0\(10),
clk => N_8,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_0_16_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI_0\(10),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_16__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_252: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.FPI.LDOP_RETO_0\,
datain => \GRLFPC2_0.FPI.LDOP_0\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_FPI_LDOP_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0000")
port map (
combout => \GRLFPC2_0.FPI.LDOP_0\,
dataf => \GRLFPC2_0.R.MK.RST\,
datae => N_81563);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_253: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO_0\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0707070505070505")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\,
dataf => N_26592,
datae => N_26591,
datad => N_26534,
datac => N_81690,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_I\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_0_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_32048_1_0,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_229\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_0_RNO_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0033003000220020")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_229\(78),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO\(53),
datac => N_28952_RETO,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO\(84),
dataa => CPI_D_INST_RETO(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_0_RNO_0_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0033003000220020")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(84),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO\(1),
datac => N_28946_RETO,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_RETO\,
dataa => CPI_D_INST_RETO(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_3_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_32340_1_0,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_3_RNO_0_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0033003000220020")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(80),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO\(55),
datac => N_28950_RETO,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO\(79),
dataa => CPI_D_INST_RETO(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A12_3_RNO_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff10")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(81),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0_4__G0_4_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0_4__G0_2_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_1_0_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_31725_1_0,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_1_0_RNO_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff10")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(81),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0_4__G0_4_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0_4__G0_2_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_1_0_RNO_0_25_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0033003000220020")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(80),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO\(55),
datac => N_28950_RETO,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO\(79),
dataa => CPI_D_INST_RETO(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_31921_1_0,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_RNO_0_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0033003000220020")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(80),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO\(55),
datac => N_28950_RETO,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO\(79),
dataa => CPI_D_INST_RETO(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_RNO_27_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff10")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(81),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0_4__G0_4_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0_4__G0_2_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_1_10_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_54_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(54),
datain => N_80636,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_22_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(22),
datain => N_80668,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_SUB_0_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffff000000ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(58),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(19),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(8));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_58_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(58),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(58),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_19_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(19),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_8_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(8),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(8),
clk => N_8,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_2_10_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_2\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_25_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(25),
datain => N_80665,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_57_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(57),
datain => N_80633,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_1_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_3_10_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_3\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1_25_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(25),
datain => N_80665,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1_57_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(57),
datain => N_80633,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_RNIJTPE_42_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_0\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_42_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(42),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_15_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_0\(15),
datain => N_81986,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2_RNILTPE_42_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_1\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2_42_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(42),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_1_15_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_1\(15),
datain => N_81986,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3_RNIOTPE_42_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_2\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3_42_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(42),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_2_15_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_2\(15),
datain => N_81986,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4_RNIQTPE_42_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_3\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4_42_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(42),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_3_15_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_3\(15),
datain => N_81986,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcfc3030fccc3000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_0\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10936_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10939_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_RNO_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0f0f00000f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_0\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M13\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM12\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_COUNTSUCCESSIVEZERO36_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datad => N_79982,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_10\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_9\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ccccff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10936_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(243));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_RNO_0_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10939_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_31_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(31),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__I0_I_0\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcfc3030fccc3000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_1\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10936_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10939_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3_RNO_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0f0f00000f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_1\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M13\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM12\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_COUNTSUCCESSIVEZERO36_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datad => N_79982,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_10\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_9\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ccccff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10936_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(243));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3_RNO_0_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10939_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_31_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(31),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__I0_I_0\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_4\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_4_10_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_4\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_53_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(53),
datain => N_80637,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_21_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(21),
datain => N_80669,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_0_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_5_10_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_5\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1_53_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(53),
datain => N_80637,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1_21_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(21),
datain => N_80669,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_1_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_6_10_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_6\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_2_53_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(53),
datain => N_80637,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_2_21_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(21),
datain => N_80669,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_7_10_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_7\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_55_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(55),
datain => N_80635,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_23_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(23),
datain => N_80667,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_0_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_8\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_8_10_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_8\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1_55_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(55),
datain => N_80635,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1_23_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(23),
datain => N_80667,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_1_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_9\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_9_10_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_9\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_2_55_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(55),
datain => N_80635,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_2_23_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(23),
datain => N_80667,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcf0fcff0c000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10944_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2_0\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(241));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0fc00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10944_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(43),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7782_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_RNO_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ffffff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2_0\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_32_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(32),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2_31_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(31),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__I0_I_0\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_241_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(241),
datain => N_36369,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcf0fcff0c000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10944_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(241));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0fc00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10944_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(43),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7782_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3_RNO_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ffffff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2_1\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_32_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(32),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3_31_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(31),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__I0_I_0\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1_241_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(241),
datain => N_36369,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5_RNIAFHI_42_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0f000fff0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_4\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5_42_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(42),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_4_15_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_4\(15),
datain => N_81986,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_43_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(43),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_43__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6_RNIDFHI_42_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0f000fff0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_6\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_5\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6_42_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_6\(42),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_5_15_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_5\(15),
datain => N_81986,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_43_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(43),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_43__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2S2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3ffc30ff0f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4534_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897_0\,
datad => \GRLFPC2_0.FPI.LDOP_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"4c4c4c44444c4444")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4534_0\,
dataf => N_26592,
datae => N_26591,
datad => N_26534,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_I\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0f0f03030f0303")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897_0\,
dataf => N_26592,
datae => N_26591,
datad => N_26534,
datac => N_81293,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\);
GRLFPC2_0_FPI_LDOP_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0000")
port map (
combout => \GRLFPC2_0.FPI.LDOP_2\,
dataf => \GRLFPC2_0.R.MK.RST\,
datae => N_81563);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_4_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(4),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_3_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(3),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SS0_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf0fc3000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4534_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897_1\,
datad => \GRLFPC2_0.FPI.LDOP_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"4c4c4c44444c4444")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4534_1\,
dataf => N_26592,
datae => N_26591,
datad => N_26534,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_I\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0f0f03030f0303")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897_1\,
dataf => N_26592,
datae => N_26591,
datad => N_26534,
datac => N_81293,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\);
GRLFPC2_0_FPI_LDOP_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0000")
port map (
combout => \GRLFPC2_0.FPI.LDOP_3\,
dataf => \GRLFPC2_0.R.MK.RST\,
datae => N_81563);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_4_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(4),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_3_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(3),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN24_ZERO_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000f33")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_0\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_0\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_3\(21),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_3\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_1_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_0\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_2_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_0\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_10_10_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_0\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_0\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_3_21_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_3\(21),
datain => N_80669,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_3_53_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_3\(53),
datain => N_80637,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN18_ZERO_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f33ffffffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_1\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_4\(21),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_4\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_2_5_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_1\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_3_6_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_1\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_11_10_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_1\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_0\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_4_21_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_4\(21),
datain => N_80669,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_4_53_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_4\(53),
datain => N_80637,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff000000ff300030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19_0\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10937_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(32),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_NORMDETECT_NOTSLFROMNORM_19_0_A2_0_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00fc00cf00ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19_0\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M13\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM12\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff00f0f0f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10937_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4_31_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(31),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__I0_I_0\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2_32_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(32),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2_43_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(43),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_43__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff000000ff300030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19_1\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10937_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(32),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_NORMDETECT_NOTSLFROMNORM_19_0_A2_1_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00fc00cf00ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19_1\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M13\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM12\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff00f0f0f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10937_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5_31_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(31),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__I0_I_0\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3_32_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(32),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3_43_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(43),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_43__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7_RNI2LRJ_42_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c0c0c0c0c0c0c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN12_SRTOSTICKY_3_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_6\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_7\(42));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN12_SRTOSTICKY: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN12_SRTOSTICKY_3_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(9),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_6_15_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_6\(15),
datain => N_81986,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7_42_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_7\(42),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333cccc0ff00ff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_12_10_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_2\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_0\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_2_25_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(25),
datain => N_80665,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_56_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(56),
datain => N_80634,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_2_57_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(57),
datain => N_80633,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_24_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(24),
datain => N_80666,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_131_RNI6FJF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00000000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10808_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G0_I_0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349_I_0_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_131: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0_0\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_RETI_0\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_254: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G0_I_0_0\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G0_I_0_RETI\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_132: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349_I_0_0\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349_I_0_RETI\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A2_RNINQ432_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff10")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(81),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_0\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_5_RNIIU4N_0_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf0fcf0fcf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2809_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_5_2_RETO\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_729_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_12_RNIJ9FU_0_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf0fcfcfefafefe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_217_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_455_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2555_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_4_0_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A2_3_0_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3cccffff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_0\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_2_RETO\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2466_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A2_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"4040404040404000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2463_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2462_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_4_0_RETO\(4),
datac => N_31763_1_RETO,
datab => N_31723_1_RETO,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_255_RETO\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A3_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffffffdf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_0\,
dataf => N_79998_RETO,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_13_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00c000c000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_1\,
datad => CPI_D_INST_RETO(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_377_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_13_C_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_13_0_RNILR152_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff10")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(81),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_5_RNIIU4N_1_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf0fcf0fcf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2809_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_5_2_RETO\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_729_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_12_RNIJ9FU_1_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf0fcfcfefafefe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_217_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_455_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2555_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_4_0_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A2_3_1_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3cccffff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_1\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_2_RETO\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2466_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A2_0_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"4040404040404000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2463_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2462_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_4_0_RETO\(4),
datac => N_31763_1_RETO,
datab => N_31723_1_RETO,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_255_RETO\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A3_0_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffffffdf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_1\,
dataf => N_79998_RETO,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_13_0_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00c000c000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_1\,
datad => CPI_D_INST_RETO(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_377_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_13_C_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_13_2_RNI3S352_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff10")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(81),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_5_RNIIU4N_9_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf0fcf0fcf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2809_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_5_2_RETO\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_729_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_12_RNIJ9FU_7_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf0fcfcfefafefe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_217_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_455_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2555_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_4_0_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A2_3_3_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3cccffff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_2\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_2_RETO\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2466_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A2_1_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"4040404040404000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2463_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2462_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_4_0_RETO\(4),
datac => N_31763_1_RETO,
datab => N_31723_1_RETO,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_255_RETO\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A3_1_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffffffdf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_2\,
dataf => N_79998_RETO,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_13_2_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00c000c000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_1\,
datad => CPI_D_INST_RETO(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_377_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_13_C_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_13_3_RNIJC652_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff10")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(81),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_3\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_5_RNIIU4N_8_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf0fcf0fcf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2809_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_5_2_RETO\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_729_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_12_RNIJ9FU_6_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf0fcfcfefafefe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_217_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_455_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2555_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_4_0_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A2_3_4_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3cccffff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_3\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_2_RETO\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2466_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A2_4_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"4040404040404000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2463_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2462_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_4_0_RETO\(4),
datac => N_31763_1_RETO,
datab => N_31723_1_RETO,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_255_RETO\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A3_2_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffffffdf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_3\,
dataf => N_79998_RETO,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_13_3_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00c000c000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_1\,
datad => CPI_D_INST_RETO(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_377_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_13_C_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_13_4_RNI0D852_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff10")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(81),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_4\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_4\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_4\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_5_RNIIU4N_7_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf0fcf0fcf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2809_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_5_2_RETO\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_729_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_12_RNIJ9FU_5_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf0fcfcfefafefe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_217_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_455_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2555_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_4_0_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A2_3_5_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3cccffff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_4\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_2_RETO\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2466_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A2_6_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"4040404040404000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2463_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2462_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_4_0_RETO\(4),
datac => N_31763_1_RETO,
datab => N_31723_1_RETO,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_255_RETO\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A3_3_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffffffdf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_4\,
dataf => N_79998_RETO,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_13_4_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00c000c000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_1\,
datad => CPI_D_INST_RETO(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_377_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_13_C_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_13_5_RNIAT952_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff10")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(81),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_5\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_5\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_5\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_5_RNIIU4N_6_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf0fcf0fcf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2809_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_5_2_RETO\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_729_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_12_RNIJ9FU_4_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf0fcfcfefafefe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_217_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_455_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2555_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_4_0_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A2_3_6_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3cccffff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_5\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_2_RETO\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2466_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A2_7_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"4040404040404000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2463_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2462_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_4_0_RETO\(4),
datac => N_31763_1_RETO,
datab => N_31723_1_RETO,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_255_RETO\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A3_4_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffffffdf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_5\,
dataf => N_79998_RETO,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_13_5_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00c000c000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_1\,
datad => CPI_D_INST_RETO(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_377_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_13_C_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_13_6_RNIQDC52_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff10")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(81),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_6\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_6\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_6\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_6\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_6\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_5_RNIIU4N_5_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf0fcf0fcf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2809_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_5_2_RETO\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_729_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_12_RNIJ9FU_3_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf0fcfcfefafefe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_217_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_455_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2555_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_4_0_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A2_3_7_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3cccffff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_6\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_2_RETO\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2466_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A2_8_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"4040404040404000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2463_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2462_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_4_0_RETO\(4),
datac => N_31763_1_RETO,
datab => N_31723_1_RETO,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_255_RETO\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A3_7_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffffffdf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_6\,
dataf => N_79998_RETO,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_13_6_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00c000c000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_1\,
datad => CPI_D_INST_RETO(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_377_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_13_C_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_13_7_RNI4UD52_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff10")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(81),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_7\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_7\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_7\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_7\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_5_RNIIU4N_4_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf0fcf0fcf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2809_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_5_2_RETO\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_729_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_12_RNIJ9FU_2_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf0fcfcfefafefe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_217_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_455_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2555_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_4_0_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A2_3_8_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3cccffff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_7\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_2_RETO\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2466_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A2_9_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"4040404040404000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2463_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2462_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_4_0_RETO\(4),
datac => N_31763_1_RETO,
datab => N_31723_1_RETO,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_255_RETO\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A3_8_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffffffdf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_7\,
dataf => N_79998_RETO,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_13_7_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00c000c000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_1\,
datad => CPI_D_INST_RETO(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_377_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_13_C_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_13_8_RNI8ON42_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff10")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(81),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_8\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_8\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_8\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_8\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_8\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_5_RNIIU4N_3_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf0fcf0fcf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2809_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_5_2_RETO\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_729_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_12_RNIK9FU_0_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf0fcfcfefafefe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_217_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_455_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2555_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_4_0_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A2_3_9_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3cccffff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_8\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_2_RETO\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2466_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A2_10_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"4040404040404000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2463_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2462_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_4_0_RETO\(4),
datac => N_31763_1_RETO,
datab => N_31723_1_RETO,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_255_RETO\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A3_9_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffffffdf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_8\,
dataf => N_79998_RETO,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_13_8_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00c000c000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_1\,
datad => CPI_D_INST_RETO(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_377_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_13_C_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A2_3_10_RNIR5P12_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff10")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(81),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_9\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_9\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_9\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_9\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_9\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_9\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_5_RNIIU4N_2_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf0fcf0fcf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_9\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2809_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_5_2_RETO\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_729_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_12_RNIK9FU_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf0fcfcfefafefe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_9\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_217_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_455_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2555_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_4_0_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A2_3_10_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3cccffff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_9\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_2_RETO\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2466_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A2_11_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"4040404040404000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_9\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2463_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2462_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_4_0_RETO\(4),
datac => N_31763_1_RETO,
datab => N_31723_1_RETO,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_255_RETO\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_A3_11_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffffffdf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_9\,
dataf => N_79998_RETO,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_I_O3_13_9_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00c000c000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_9\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_1\,
datad => CPI_D_INST_RETO(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_377_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O3_13_C_RETO\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_RNI4COD1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(84),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_0\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_0\,
datac => N_28946_RETO_0,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_RETO_0\,
dataa => CPI_D_INST_RETO_0(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_22_RNIGNLN_7: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_0\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_RETO\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_133: stratixii_lcell_ff port map (
regout => N_28946_RETO_0,
datain => N_28946,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_134: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_RETO_0\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_135: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_0(9),
datain => N_59,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_136_RNIO7QG1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(84),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_1\,
datac => N_28946_RETO_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_RETO_1\,
dataa => CPI_D_INST_RETO_1(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_22_RNIGNLN_6: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_1\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_RETO\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_136: stratixii_lcell_ff port map (
regout => N_28946_RETO_1,
datain => N_28946,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_137: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_RETO_1\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_138: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_1(9),
datain => N_59,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_139_RNIHFQG1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(84),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_2\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_2\,
datac => N_28946_RETO_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_RETO_2\,
dataa => CPI_D_INST_RETO_2(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_22_RNIGNLN_5: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_2\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_RETO\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_139: stratixii_lcell_ff port map (
regout => N_28946_RETO_2,
datain => N_28946,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_140: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_RETO_2\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_141: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_2(9),
datain => N_59,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_142_RNIKJQG1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(84),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_3\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_3\,
datac => N_28946_RETO_3,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_RETO_3\,
dataa => CPI_D_INST_RETO_3(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_22_RNIGNLN_4: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_3\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_RETO\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_142: stratixii_lcell_ff port map (
regout => N_28946_RETO_3,
datain => N_28946,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_143: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_RETO_3\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_144: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_3(9),
datain => N_59,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_145_RNIVJQG1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(84),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_4\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_4\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_4\,
datac => N_28946_RETO_4,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_RETO_4\,
dataa => CPI_D_INST_RETO_4(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_4: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_4: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_22_RNIGNLN_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_4\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_RETO\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_145: stratixii_lcell_ff port map (
regout => N_28946_RETO_4,
datain => N_28946,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_146: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_RETO_4\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_147: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_4(9),
datain => N_59,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_148_RNI1OQG1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(84),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_5\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_5\,
datac => N_28946_RETO_5,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_RETO_5\,
dataa => CPI_D_INST_RETO_5(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_5: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_5: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_22_RNIGNLN_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_5\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_RETO\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_148: stratixii_lcell_ff port map (
regout => N_28946_RETO_5,
datain => N_28946,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_149: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_RETO_5\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_150: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_5(9),
datain => N_59,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_151_RNIQVQG1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(84),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_6\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_6\,
datac => N_28946_RETO_6,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_RETO_6\,
dataa => CPI_D_INST_RETO_6(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_6: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_6: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_22_RNIGNLN_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_6\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_RETO\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_151: stratixii_lcell_ff port map (
regout => N_28946_RETO_6,
datain => N_28946,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_152: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_RETO_6\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_153: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_6(9),
datain => N_59,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_154_RNI50RG1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(84),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_7\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_7\,
datac => N_28946_RETO_7,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_RETO_7\,
dataa => CPI_D_INST_RETO_7(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_7: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_7: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_22_RNIGNLN_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_7\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_RETO\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_154: stratixii_lcell_ff port map (
regout => N_28946_RETO_7,
datain => N_28946,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_155: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_RETO_7\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_156: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_7(9),
datain => N_59,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_157_RNIKI1D2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff003caabe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(82),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_8\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(82),
dataa => CPI_D_INST_RETO_0(11));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_12_RNIK9SJ1_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000fffc0200fefc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(65),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_8: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_8: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_157: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO_0\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_158: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(82),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_159: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_0(11),
datain => N_61,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_160_RNI4U1D2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff003caabe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(82),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_9\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_9\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(82),
dataa => CPI_D_INST_RETO_1(11));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_12_RNIK9SJ1_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000fffc0200fefc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(65),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_9: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_9\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_9: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_9\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_160: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO_1\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_161: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(82),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_162: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_1(11),
datain => N_61,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_10_RNI9L672: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff003caabe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(82),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_10\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_10\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_2\(82),
dataa => CPI_D_INST_RETO_2(11));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_12_RNIK9SJ1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000fffc0200fefc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(65),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_10: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_10\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_10: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_10\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_163: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO_2\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_164: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_2\(82),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_165: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_2(11),
datain => N_61,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_11_RNIKL672: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff003caabe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(82),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO_3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_11\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_11\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_3\(82),
dataa => CPI_D_INST_RETO_3(11));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_12_RNIK9SJ1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000fffc0200fefc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(65),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_11: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_11\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_11: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_11\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_166: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO_3\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_167: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_3\(82),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_168: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_3(11),
datain => N_61,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_12_RNIDT672: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff003caabe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(82),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO_4\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_12\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_12\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO_4\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_4\(82),
dataa => CPI_D_INST_RETO_4(11));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_12_RNIK9SJ1_7: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000fffc0200fefc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(65),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_12: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_12\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_12: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_12\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_169: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO_4\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_170: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_4\(82),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_171: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_4(11),
datain => N_61,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_13_RNIF1772: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff003caabe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(82),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_13\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_13\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO_5\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_5\(82),
dataa => CPI_D_INST_RETO_5(11));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_12_RNIK9SJ1_6: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000fffc0200fefc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(65),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_13: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_13\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_13: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_13\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_172: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO_5\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_173: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_5\(82),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_174: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_5(11),
datain => N_61,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_14_RNIQ1772: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff003caabe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(82),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_14\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_14\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO_6\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_6\(82),
dataa => CPI_D_INST_RETO_6(11));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_12_RNIK9SJ1_5: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000fffc0200fefc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(65),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_14: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_14\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_14: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_14\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_175: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO_6\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_176: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_6\(82),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_177: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_6(11),
datain => N_61,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_15_RNIS5772: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff003caabe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_157\(82),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_15\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_15\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO_7\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_7\(82),
dataa => CPI_D_INST_RETO_7(11));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_12_RNIK9SJ1_4: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000fffc0200fefc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(65),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_15: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_15\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_15: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_15\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_178: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO_7\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_179: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_7\(82),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_180: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_7(11),
datain => N_61,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_16_RNILD772: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff003caabe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_158\(82),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO_8\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_16\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_16\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO_8\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_8\(82),
dataa => CPI_D_INST_RETO_8(11));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_12_RNIK9SJ1_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000fffc0200fefc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(65),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_16: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_16\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_16: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_16\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_181: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2_RETO_8\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO2\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_182: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_8\(82),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_183: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_8(11),
datain => N_61,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_17_RNIHGFL2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f0c0a08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_147\(83),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_0\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_17\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_17\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_0\(2),
datab => N_28947_RETO_0,
dataa => CPI_D_INST_RETO_0(7));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_17: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_17\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_17: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_17\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_26_RNI5C422_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000fa0033")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_0\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_I_0_0_RETO\,
datac => \GRLFPC2_0.FPO.FRAC_RETO\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0_RETO\(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_184: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_0\(2),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M\(2),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_185: stratixii_lcell_ff port map (
regout => N_28947_RETO_0,
datain => N_28947,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_186: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_0(7),
datain => N_57,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_18_RNISGFL2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f0c0a08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_148\(83),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_1\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_18\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_18\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_1\(2),
datab => N_28947_RETO_1,
dataa => CPI_D_INST_RETO_1(7));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_18: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_18\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_18: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_18\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_26_RNI5C422: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000fa0033")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_1\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_I_0_0_RETO\,
datac => \GRLFPC2_0.FPO.FRAC_RETO\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0_RETO\(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_187: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_1\(2),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M\(2),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_188: stratixii_lcell_ff port map (
regout => N_28947_RETO_1,
datain => N_28947,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_189: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_1(7),
datain => N_57,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_19_RNI6VDL2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f0c0a08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_149\(83),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_2\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_19\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_19\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_2\(2),
datab => N_28947_RETO_2,
dataa => CPI_D_INST_RETO_2(7));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_19: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_19\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_19: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_19\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_26_RNIVE222_6: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000fa0033")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_2\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_I_0_0_RETO\,
datac => \GRLFPC2_0.FPO.FRAC_RETO\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0_RETO\(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_190: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_2\(2),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M\(2),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_191: stratixii_lcell_ff port map (
regout => N_28947_RETO_2,
datain => N_28947,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_192: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_2(7),
datain => N_57,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_20_RNIV2EL2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f0c0a08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_150\(83),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_3\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_20\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_20\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_3\(2),
datab => N_28947_RETO_3,
dataa => CPI_D_INST_RETO_3(7));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_20: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_20\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_20: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_20\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_26_RNIVE222_5: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000fa0033")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_3\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_I_0_0_RETO\,
datac => \GRLFPC2_0.FPO.FRAC_RETO\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0_RETO\(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_193: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_3\(2),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M\(2),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_194: stratixii_lcell_ff port map (
regout => N_28947_RETO_3,
datain => N_28947,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_195: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_3(7),
datain => N_57,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_21_RNIA3EL2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f0c0a08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_151\(83),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_4\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_21\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_21\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_4\(2),
datab => N_28947_RETO_4,
dataa => CPI_D_INST_RETO_4(7));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_21: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_21\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_21: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_21\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_26_RNIVE222_4: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000fa0033")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_4\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_I_0_0_RETO\,
datac => \GRLFPC2_0.FPO.FRAC_RETO\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0_RETO\(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_196: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_4\(2),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M\(2),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_197: stratixii_lcell_ff port map (
regout => N_28947_RETO_4,
datain => N_28947,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_198: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_4(7),
datain => N_57,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_22_RNIHQBL2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f0c0a08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_152\(83),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_5\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_22\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_22\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_5\(2),
datab => N_28947_RETO_5,
dataa => CPI_D_INST_RETO_5(7));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_22: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_22\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_22: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_22\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_26_RNIVE222_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000fa0033")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_5\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_I_0_0_RETO\,
datac => \GRLFPC2_0.FPO.FRAC_RETO\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0_RETO\(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_199: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_5\(2),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M\(2),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_200: stratixii_lcell_ff port map (
regout => N_28947_RETO_5,
datain => N_28947,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_201: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_5(7),
datain => N_57,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_23_RNIAMAL2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f0c0a08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_153\(83),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_6\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_23\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_23\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_6\(2),
datab => N_28947_RETO_6,
dataa => CPI_D_INST_RETO_6(7));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_23: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_23\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_23: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_23\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_26_RNIVE222_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000fa0033")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_6\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_I_0_0_RETO\,
datac => \GRLFPC2_0.FPO.FRAC_RETO\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0_RETO\(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_202: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_6\(2),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M\(2),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_203: stratixii_lcell_ff port map (
regout => N_28947_RETO_6,
datain => N_28947,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_204: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_6(7),
datain => N_57,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_24_RNILMAL2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f0c0a08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_154\(83),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_7\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_24\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_24\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_7\(2),
datab => N_28947_RETO_7,
dataa => CPI_D_INST_RETO_7(7));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_24: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_24\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_24: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_24\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_26_RNIVE222_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000fa0033")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_7\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_I_0_0_RETO\,
datac => \GRLFPC2_0.FPO.FRAC_RETO\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0_RETO\(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_205: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_7\(2),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M\(2),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_206: stratixii_lcell_ff port map (
regout => N_28947_RETO_7,
datain => N_28947,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_207: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_7(7),
datain => N_57,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_25_RNINQAL2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f0c0a08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_155\(83),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_8\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_25\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_25\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_8\(2),
datab => N_28947_RETO_8,
dataa => CPI_D_INST_RETO_8(7));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_25: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_25\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_25: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_25\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_26_RNIVE222_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000fa0033")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_8\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_I_0_0_RETO\,
datac => \GRLFPC2_0.FPO.FRAC_RETO\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0_RETO\(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_208: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_8\(2),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M\(2),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_209: stratixii_lcell_ff port map (
regout => N_28947_RETO_8,
datain => N_28947,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_210: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_8(7),
datain => N_57,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_26_RNIG2BL2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f0c0a08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_156\(83),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_9\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_26\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_26\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_9\(2),
datab => N_28947_RETO_9,
dataa => CPI_D_INST_RETO_9(7));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_26: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_26\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_26: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_26\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_26_RNIVE222: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000fa0033")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_9\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_I_0_0_RETO\,
datac => \GRLFPC2_0.FPO.FRAC_RETO\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0_RETO\(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_211: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_9\(2),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M\(2),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_212: stratixii_lcell_ff port map (
regout => N_28947_RETO_9,
datain => N_28947,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_213: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_9(7),
datain => N_57,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_27_RNIT3TH2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f0c0a08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_280\(85),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_27\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_27\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO_0\,
datab => N_28945_RETO_0,
dataa => CPI_D_INST_RETO_0(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_1_RNI1GKU1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000dd000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_0\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_I_0_0_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_RETO\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5330_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_27: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_27\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_27: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_27\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_214: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO_0\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_215: stratixii_lcell_ff port map (
regout => N_28945_RETO_0,
datain => N_28945,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_216: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_0(10),
datain => N_60,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_28_RNI84TH2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f0c0a08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_281\(85),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_28\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_28\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO_1\,
datab => N_28945_RETO_1,
dataa => CPI_D_INST_RETO_1(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_1_RNI1GKU1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000dd000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_1\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_I_0_0_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_RETO\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5330_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_28: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_28\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_28: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_28\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_217: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO_1\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_218: stratixii_lcell_ff port map (
regout => N_28945_RETO_1,
datain => N_28945,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_219: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_1(10),
datain => N_60,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_29_RNIIIRH2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f0c0a08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_282\(85),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_2\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_29\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_29\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO_2\,
datab => N_28945_RETO_2,
dataa => CPI_D_INST_RETO_2(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_1_RNIRIIU1_5: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000dd000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_2\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_I_0_0_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_RETO\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5330_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_29: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_29\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_29: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_29\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_220: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO_2\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_221: stratixii_lcell_ff port map (
regout => N_28945_RETO_2,
datain => N_28945,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_222: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_2(10),
datain => N_60,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_30_RNIBMRH2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f0c0a08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_283\(85),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_3\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_30\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_30\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO_3\,
datab => N_28945_RETO_3,
dataa => CPI_D_INST_RETO_3(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_1_RNIRIIU1_4: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000dd000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_3\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_I_0_0_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_RETO\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5330_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_30: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_30\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_30: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_30\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_223: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO_3\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_224: stratixii_lcell_ff port map (
regout => N_28945_RETO_3,
datain => N_28945,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_225: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_3(10),
datain => N_60,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_31_RNIMMRH2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f0c0a08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_284\(85),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_4\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_31\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_31\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO_4\,
datab => N_28945_RETO_4,
dataa => CPI_D_INST_RETO_4(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_1_RNIRIIU1_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000dd000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_4\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_I_0_0_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_RETO\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5330_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_31: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_31\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_31: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_31\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_226: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO_4\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_227: stratixii_lcell_ff port map (
regout => N_28945_RETO_4,
datain => N_28945,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_228: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_4(10),
datain => N_60,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_32_RNIFURH2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f0c0a08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_285\(85),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_5\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_32\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_32\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO_5\,
datab => N_28945_RETO_5,
dataa => CPI_D_INST_RETO_5(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_1_RNIRIIU1_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000dd000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_5\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_I_0_0_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_RETO\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5330_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_32: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_32\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_32: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_32\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_229: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO_5\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_230: stratixii_lcell_ff port map (
regout => N_28945_RETO_5,
datain => N_28945,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_231: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_5(10),
datain => N_60,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_33_RNIH2SH2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f0c0a08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_286\(85),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_6\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_33\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_33\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO_6\,
datab => N_28945_RETO_6,
dataa => CPI_D_INST_RETO_6(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_1_RNIRIIU1_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000dd000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_6\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_I_0_0_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_RETO\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5330_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_33: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_33\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_33: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_33\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_232: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO_6\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_233: stratixii_lcell_ff port map (
regout => N_28945_RETO_6,
datain => N_28945,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_234: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_6(10),
datain => N_60,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_34_RNIS2SH2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f0c0a08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_287\(85),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_7\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_34\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_34\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO_7\,
datab => N_28945_RETO_7,
dataa => CPI_D_INST_RETO_7(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_1_RNIRIIU1_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000dd000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_7\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_I_0_0_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_RETO\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5330_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_34: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_34\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_34: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_34\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_235: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO_7\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_236: stratixii_lcell_ff port map (
regout => N_28945_RETO_7,
datain => N_28945,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_237: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_7(10),
datain => N_60,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_35_RNIU6SH2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f0c0a08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_288\(85),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_8\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_35\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_35\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO_8\,
datab => N_28945_RETO_8,
dataa => CPI_D_INST_RETO_8(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_1_RNIRIIU1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000dd000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO_8\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_I_0_0_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_RETO\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5330_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_35: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_35\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_35: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_35\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_238: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_RETO_8\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_239: stratixii_lcell_ff port map (
regout => N_28945_RETO_8,
datain => N_28945,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_240: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_8(10),
datain => N_60,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_36_RNIGNVA1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(80),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_36\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_0\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_36\,
datac => N_28950_RETO_0,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO_0\(79),
dataa => CPI_D_INST_RETO_0(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_36: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_36\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_36: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_36\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_79_RNIKRLN_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_0\(55),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_241: stratixii_lcell_ff port map (
regout => N_28950_RETO_0,
datain => N_28950,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_242: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO_0\(79),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M\(79),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_243: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_0(5),
datain => N_55,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_37_RNIRNVA1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(80),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_37\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_1\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_37\,
datac => N_28950_RETO_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO_1\(79),
dataa => CPI_D_INST_RETO_1(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_37: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_37\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_37: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_37\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_79_RNIKRLN_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_1\(55),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_244: stratixii_lcell_ff port map (
regout => N_28950_RETO_1,
datain => N_28950,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_245: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO_1\(79),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M\(79),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_246: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_1(5),
datain => N_55,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_38_RNIQMHE1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_38\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_2\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_38\,
datac => N_28950_RETO_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO_2\(79),
dataa => CPI_D_INST_RETO_2(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_38: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_38\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_38: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_38\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_79_RNI8Q7R_4: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_2\(55),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_247: stratixii_lcell_ff port map (
regout => N_28950_RETO_2,
datain => N_28950,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_248: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO_2\(79),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M\(79),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_249: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_2(5),
datain => N_55,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_39_RNIA2IE1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_39\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_3\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_39\,
datac => N_28950_RETO_3,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO_3\(79),
dataa => CPI_D_INST_RETO_3(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_39: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bbabffffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_39\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_39: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_39\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_79_RNI8Q7R_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_3\(55),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_250: stratixii_lcell_ff port map (
regout => N_28950_RETO_3,
datain => N_28950,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_251: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO_3\(79),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M\(79),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_252: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_3(5),
datain => N_55,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_40_RNI36IE1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_40\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_4\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_40\,
datac => N_28950_RETO_4,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO_4\(79),
dataa => CPI_D_INST_RETO_4(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_40: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"afabffffafafffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_40\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_40: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_40\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_79_RNI8Q7R_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_4\(55),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_253: stratixii_lcell_ff port map (
regout => N_28950_RETO_4,
datain => N_28950,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_254: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO_4\(79),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M\(79),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_255: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_4(5),
datain => N_55,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_41_RNIE6IE1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_41\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_5\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_41\,
datac => N_28950_RETO_5,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO_5\(79),
dataa => CPI_D_INST_RETO_5(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_41: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"afabffffafafffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_41\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_41: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_41\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_79_RNI8Q7R_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_5\(55),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_256: stratixii_lcell_ff port map (
regout => N_28950_RETO_5,
datain => N_28950,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_257: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO_5\(79),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M\(79),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_258: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_5(5),
datain => N_55,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_42_RNI7EIE1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_42\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_6\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_42\,
datac => N_28950_RETO_6,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO_6\(79),
dataa => CPI_D_INST_RETO_6(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_42: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"afabffffafafffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_42\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_42: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_42\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_79_RNI8Q7R_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_6\(55),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_259: stratixii_lcell_ff port map (
regout => N_28950_RETO_6,
datain => N_28950,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_260: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO_6\(79),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M\(79),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_261: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_6(5),
datain => N_55,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_43_RNI9IIE1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_43\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_7\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_43\,
datac => N_28950_RETO_7,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO_7\(79),
dataa => CPI_D_INST_RETO_7(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_43: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"afabffffafafffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_43\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_43: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_43\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_79_RNI8Q7R: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_7\(55),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_262: stratixii_lcell_ff port map (
regout => N_28950_RETO_7,
datain => N_28950,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_263: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO_7\(79),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M\(79),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_264: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_7(5),
datain => N_55,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_44_RNILIIE1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_44\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_8\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_44\,
datac => N_28950_RETO_8,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO_8\(79),
dataa => CPI_D_INST_RETO_8(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_44: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"afabffffafafffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_44\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_44: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_44\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_79_RNI9Q7R: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_8\(55),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_265: stratixii_lcell_ff port map (
regout => N_28950_RETO_8,
datain => N_28950,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_266: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO_8\(79),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M\(79),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_267: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_8(5),
datain => N_55,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_45_RNITN0B1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(79),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_45\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_0\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_45\,
datac => N_28951_RETO_0,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_0\(6),
dataa => CPI_D_INST_RETO_0(8));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_45: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"afabffffafafffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_45\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_45: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_45\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_38_RNIFRLN_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_0\(54),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_268: stratixii_lcell_ff port map (
regout => N_28951_RETO_0,
datain => N_28951,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_269: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_0\(6),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M\(6),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_270: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_0(8),
datain => N_58,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_46_RNIMV0B1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_245\(79),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_46\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_1\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_46\,
datac => N_28951_RETO_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_1\(6),
dataa => CPI_D_INST_RETO_1(8));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_46: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"afabffffafafffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_46\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_46: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_46\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_38_RNIFRLN: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_1\(54),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_271: stratixii_lcell_ff port map (
regout => N_28951_RETO_1,
datain => N_28951,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_272: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_1\(6),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M\(6),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_273: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_1(8),
datain => N_58,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_47_RNILUIE1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_246\(79),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_47\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_2\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_47\,
datac => N_28951_RETO_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_2\(6),
dataa => CPI_D_INST_RETO_2(8));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_47: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"afabffffafafffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_47\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_47: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_47\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_38_RNI3Q7R_4: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_2\(54),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_274: stratixii_lcell_ff port map (
regout => N_28951_RETO_2,
datain => N_28951,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_275: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_2\(6),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M\(6),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_276: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_2(8),
datain => N_58,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_48_RNI0VIE1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_247\(79),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_48\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_3\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_48\,
datac => N_28951_RETO_3,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_3\(6),
dataa => CPI_D_INST_RETO_3(8));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_48: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"afabffffafafffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_48\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_48: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_48\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_38_RNI3Q7R_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_3\(54),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_277: stratixii_lcell_ff port map (
regout => N_28951_RETO_3,
datain => N_28951,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_278: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_3\(6),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M\(6),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_279: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_3(8),
datain => N_58,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_49_RNIGAJE1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(79),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_49\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_4\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_49\,
datac => N_28951_RETO_4,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_4\(6),
dataa => CPI_D_INST_RETO_4(8));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_49: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"afabffffafafffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_49\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_49: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_49\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_38_RNI3Q7R_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_4\(54),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_280: stratixii_lcell_ff port map (
regout => N_28951_RETO_4,
datain => N_28951,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_281: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_4\(6),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M\(6),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_282: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_4(8),
datain => N_58,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_50_RNI9EJE1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(79),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_50\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_5\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_50\,
datac => N_28951_RETO_5,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_5\(6),
dataa => CPI_D_INST_RETO_5(8));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_50: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"afabffffafafffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_50\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_50: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_50\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_38_RNI3Q7R_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_5\(54),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_283: stratixii_lcell_ff port map (
regout => N_28951_RETO_5,
datain => N_28951,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_284: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_5\(6),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M\(6),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_285: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_5(8),
datain => N_58,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_51_RNIKEJE1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(79),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_51\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_6\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_51\,
datac => N_28951_RETO_6,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_6\(6),
dataa => CPI_D_INST_RETO_6(8));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_51: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"afabffffafafffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_51\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_51: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_51\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_38_RNI3Q7R_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_6\(54),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_286: stratixii_lcell_ff port map (
regout => N_28951_RETO_6,
datain => N_28951,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_287: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_6\(6),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M\(6),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_288: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_6(8),
datain => N_58,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_52_RNIDMJE1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_52\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_7\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_52\,
datac => N_28951_RETO_7,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_7\(6),
dataa => CPI_D_INST_RETO_7(8));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_52: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"afabffffafafffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_52\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_52: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_52\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_38_RNI3Q7R: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_7\(54),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_289: stratixii_lcell_ff port map (
regout => N_28951_RETO_7,
datain => N_28951,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_290: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_7\(6),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M\(6),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_291: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_7(8),
datain => N_58,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_53_RNIGQJE1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_53\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_8\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_53\,
datac => N_28951_RETO_8,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_8\(6),
dataa => CPI_D_INST_RETO_8(8));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_53: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"afabffffafafffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_53\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_53: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_53\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_38_RNI4Q7R: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_8\(54),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_292: stratixii_lcell_ff port map (
regout => N_28951_RETO_8,
datain => N_28951,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_293: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO_8\(6),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M\(6),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_294: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_8(8),
datain => N_58,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_54_RNIAS1B1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_230\(78),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_54\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_0\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_54\,
datac => N_28952_RETO_0,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO_0\(84),
dataa => CPI_D_INST_RETO_0(12));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_54: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"afabffffafafffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_54\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_54: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_54\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_78_RNIJRLN_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_0\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_295: stratixii_lcell_ff port map (
regout => N_28952_RETO_0,
datain => N_28952,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_296: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO_0\(84),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M\(84),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_297: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_0(12),
datain => N_62,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_55_RNI3O0B1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_231\(78),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_55\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_1\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_55\,
datac => N_28952_RETO_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO_1\(84),
dataa => CPI_D_INST_RETO_1(12));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_55: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"afabffffafafffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_55\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_55: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_55\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_78_RNIJRLN_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_1\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_298: stratixii_lcell_ff port map (
regout => N_28952_RETO_1,
datain => N_28952,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_299: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO_1\(84),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M\(84),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_300: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_1(12),
datain => N_62,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_56_RNIAFUA1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_232\(78),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_56\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_2\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_56\,
datac => N_28952_RETO_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO_2\(84),
dataa => CPI_D_INST_RETO_2(12));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_56: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"afabffffafafffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_56\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_56: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_56\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_78_RNIJRLN_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_2\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_301: stratixii_lcell_ff port map (
regout => N_28952_RETO_2,
datain => N_28952,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_302: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO_2\(84),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M\(84),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_303: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_2(12),
datain => N_62,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_57_RNI9EGE1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_233\(78),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_57\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_3\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_57\,
datac => N_28952_RETO_3,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO_3\(84),
dataa => CPI_D_INST_RETO_3(12));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_57: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"afabffffafafffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_57\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_57: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_57\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_78_RNI7Q7R_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_3\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_304: stratixii_lcell_ff port map (
regout => N_28952_RETO_3,
datain => N_28952,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_305: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO_3\(84),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M\(84),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_306: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_3(12),
datain => N_62,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_58_RNIKEGE1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_234\(78),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_58\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_4\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_58\,
datac => N_28952_RETO_4,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO_4\(84),
dataa => CPI_D_INST_RETO_4(12));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_58: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"afabffffafafffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_58\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_58: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_58\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_78_RNI7Q7R_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_4\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_307: stratixii_lcell_ff port map (
regout => N_28952_RETO_4,
datain => N_28952,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_308: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO_4\(84),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M\(84),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_309: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_4(12),
datain => N_62,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_59_RNI4QGE1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(78),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_59\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_5\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_59\,
datac => N_28952_RETO_5,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO_5\(84),
dataa => CPI_D_INST_RETO_5(12));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_59: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"afabffffafafffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_59\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_59: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_59\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_78_RNI7Q7R_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_5\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_310: stratixii_lcell_ff port map (
regout => N_28952_RETO_5,
datain => N_28952,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_311: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO_5\(84),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M\(84),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_312: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_5(12),
datain => N_62,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_60_RNITTGE1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(78),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_60\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_6\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_60\,
datac => N_28952_RETO_6,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO_6\(84),
dataa => CPI_D_INST_RETO_6(12));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_60: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"afabffffafafffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_60\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_60: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_60\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_78_RNI7Q7R_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_6\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_313: stratixii_lcell_ff port map (
regout => N_28952_RETO_6,
datain => N_28952,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_314: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO_6\(84),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M\(84),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_315: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_6(12),
datain => N_62,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_61_RNI8UGE1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(78),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_61\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_7\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_61\,
datac => N_28952_RETO_7,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO_7\(84),
dataa => CPI_D_INST_RETO_7(12));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_61: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"afabffffafafffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_61\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_61: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_61\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_78_RNI7Q7R: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_7\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_316: stratixii_lcell_ff port map (
regout => N_28952_RETO_7,
datain => N_28952,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_317: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO_7\(84),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M\(84),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_318: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_7(12),
datain => N_62,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_62_RNI26HE1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(78),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_62\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_8\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_62\,
datac => N_28952_RETO_8,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO_8\(84),
dataa => CPI_D_INST_RETO_8(12));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_0_62: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"afabffffafafffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_62\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_62: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0fff00ff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_62\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_78_RNI8Q7R: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_8\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10930_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_319: stratixii_lcell_ff port map (
regout => N_28952_RETO_8,
datain => N_28952,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_320: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M_RETO_8\(84),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_24_M\(84),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_321: stratixii_lcell_ff port map (
regout => CPI_D_INST_RETO_8(12),
datain => N_62,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN5_ZERO_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"77770fffeeeefff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_0\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_3\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_3\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_2_8_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_0\(8),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_13_10_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_3\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_0\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_3_55_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_3\(55),
datain => N_80635,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1_56_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(56),
datain => N_80634,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1_24_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(24),
datain => N_80666,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_3_23_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_3\(23),
datain => N_80667,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0c0c04040c0404")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_0\,
dataf => N_26592,
datae => N_26591,
datad => N_26534,
datac => N_81248_0,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_SUB_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000100010001")
port map (
combout => N_81248_0,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\,
datad => \GRLFPC2_0.FPI.LDOP_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff3000ffff3300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748\,
datae => \GRLFPC2_0.FPI.LDOP_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_237\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_0_68_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506_0\,
dataf => \GRLFPC2_0.FPI.LDOP_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(12),
datad => \GRLFPC2_0.R.MK.RST2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(47),
datab => N_7);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_4: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0c0c04040c0404")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118_1\,
dataf => N_26592,
datae => N_26591,
datad => N_26534,
datac => N_81248_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_SUB_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000100010001")
port map (
combout => N_81248_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\,
datad => \GRLFPC2_0.FPI.LDOP_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff3000ffff3300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748\,
datae => \GRLFPC2_0.FPI.LDOP_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_237\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_1_68_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506_1\,
dataf => \GRLFPC2_0.FPI.LDOP_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(12),
datad => \GRLFPC2_0.R.MK.RST2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(47),
datab => N_7);
GRLFPC2_0_FPI_LDOP_4: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0000")
port map (
combout => \GRLFPC2_0.FPI.LDOP_4\,
dataf => N_81563_0,
datae => \GRLFPC2_0.R.MK.RST_0\);
GRLFPC2_0_FPI_LDOP_SUB_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffdfff55ff55ff55")
port map (
combout => N_81563_0,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7612_I_A7_10\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7612_I_A7_6\,
datad => \GRLFPC2_0.R.MK.RST2\,
datac => \GRLFPC2_0.R.STATE_O_3\(0),
datab => \GRLFPC2_0.R.STATE_O_3\(1),
dataa => N_7);
GRLFPC2_0_FPI_LDOP_4_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000000000000000")
port map (
combout => \GRLFPC2_0.R.MK.RST_0\,
dataf => \GRLFPC2_0.FPO.BUSY_O\,
datae => \GRLFPC2_0.R.MK.RST_4\,
datad => \GRLFPC2_0.HOLDN_O\,
datac => \GRLFPC2_0.R.MK.HOLDN2_O\);
GRLFPC2_0_FPI_LDOP_5: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0000")
port map (
combout => \GRLFPC2_0.FPI.LDOP_5\,
dataf => N_81563_1,
datae => \GRLFPC2_0.R.MK.RST_1\);
GRLFPC2_0_FPI_LDOP_SUB_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffdfff55ff55ff55")
port map (
combout => N_81563_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7612_I_A7_10\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7612_I_A7_6\,
datad => \GRLFPC2_0.R.MK.RST2\,
datac => \GRLFPC2_0.R.STATE_O_3\(0),
datab => \GRLFPC2_0.R.STATE_O_3\(1),
dataa => N_7);
GRLFPC2_0_FPI_LDOP_5_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000000000000000")
port map (
combout => \GRLFPC2_0.R.MK.RST_1\,
dataf => \GRLFPC2_0.FPO.BUSY_O\,
datae => \GRLFPC2_0.R.MK.RST_4\,
datad => \GRLFPC2_0.HOLDN_O\,
datac => \GRLFPC2_0.R.MK.HOLDN2_O\);
GRLFPC2_0_FPI_LDOP_6: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0000")
port map (
combout => \GRLFPC2_0.FPI.LDOP_6\,
dataf => N_81563_2,
datae => \GRLFPC2_0.R.MK.RST_2\);
GRLFPC2_0_FPI_LDOP_SUB_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffdfff55ff55ff55")
port map (
combout => N_81563_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7612_I_A7_10\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7612_I_A7_6\,
datad => \GRLFPC2_0.R.MK.RST2\,
datac => \GRLFPC2_0.R.STATE_O_3\(0),
datab => \GRLFPC2_0.R.STATE_O_3\(1),
dataa => N_7);
GRLFPC2_0_FPI_LDOP_6_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000000000000000")
port map (
combout => \GRLFPC2_0.R.MK.RST_2\,
dataf => \GRLFPC2_0.FPO.BUSY_O\,
datae => \GRLFPC2_0.R.MK.RST_4\,
datad => \GRLFPC2_0.HOLDN_O\,
datac => \GRLFPC2_0.R.MK.HOLDN2_O\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_0\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_RNO_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff80")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_3\,
datad => N_33355,
datac => N_32344_1,
datab => N_27297_1,
dataa => N_31941_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_1\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_RNO_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff80")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_3\,
datad => N_33355,
datac => N_32344_1,
datab => N_27297_1,
dataa => N_31941_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2_0_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_4\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2_RNO_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff80")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_3\,
datad => N_33355,
datac => N_32344_1,
datab => N_27297_1,
dataa => N_31941_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3_0_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_5\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3_RNO_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff80")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_3\,
datad => N_33355,
datac => N_32344_1,
datab => N_27297_1,
dataa => N_31941_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4_0_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_6\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4_RNO_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff80")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_3\,
datad => N_33355,
datac => N_32344_1,
datab => N_27297_1,
dataa => N_31941_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5_0_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(0),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_8\,
clk => N_8,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5_RNO_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff80")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_3\,
datad => N_33355,
datac => N_32344_1,
datab => N_27297_1,
dataa => N_31941_1);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_322: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_0\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_0\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccc0ccc0ccc00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_647\,
datae => N_32136_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_329\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2757\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_323: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_RETO_1\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_1\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_I_0_A2_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccc0ccc0ccc00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1916_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_647\,
datae => N_32136_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_329\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2757\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_324: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(73),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3729_I_0_0\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_324_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"030303030303030f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3729_I_0_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_318\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O2_2\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O2_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(66));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_325: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(73),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3729_I_0_1\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_325_RNO: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"030303030303030f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3729_I_0_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_318\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O2_2\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_O2_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(66));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_326: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_0\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_0\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffcccf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2477\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O2_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2765\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_327: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_RETO_1\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_1\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffcccf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_2_2_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2477\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O2_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2765\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_328: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_0\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_0\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000f000f333f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_237\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_329\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_329: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_RETO_1\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_1\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000f000f333f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_0_O2_0_O3_0_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_237\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_329\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_330: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(65),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(65),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_65_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(65),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1780_I\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_331: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(65),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(65),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_65_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(65),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1780_I\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_332: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_0\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_0\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTABORTNULLEXC_0_O2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ffff00ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(76));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_333: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_1\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_1\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTABORTNULLEXC_0_O2_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ffff00ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(76));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_334: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_RETO_2\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_2\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTABORTNULLEXC_0_O2_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ffff00ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1742_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(76));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_335: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_0\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_0\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_O3_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0fff0f0cffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN11_WQSTSETS\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_336: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_1\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_1\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_O3_0_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0fff0f0cffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN11_WQSTSETS\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_337: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_RETO_2\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_2\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_O3_1_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0fff0f0cffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN11_WQSTSETS\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_338: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_RETO_0\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_0\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_UN10_SELECTEDMIPTR_I_0_O2_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff0fffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_642_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_422\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(76));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_339: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_0\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_A3_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cccccccc000ccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2807\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5065\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_6\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3848\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(46));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_340: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_1\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_1\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_A3_1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cccccccc000ccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2807\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5065\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_6\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3848\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(46));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_341: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_2\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_2\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_A3_2: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cccccccc000ccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2807\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5065\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_6\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3848\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(46));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_342: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_3\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_3\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_A3_3: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cccccccc000ccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2807\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5065\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_6\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3848\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(46));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_343: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_4\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_4\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_A3_4: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cccccccc000ccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2807\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5065\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_6\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3848\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(46));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_344: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_5\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_5\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_A3_5: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cccccccc000ccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2807\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5065\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_6\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3848\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_32141_1_0,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238_0\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251_0\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_RNO_0_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000333000002220")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251_0\(80),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5_RETO_36\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_I_M_RETO_0\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2810_RETO_36\,
datac => N_28950_RETO_0,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO_0\(79),
dataa => CPI_D_INST_RETO_0(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_RNO_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff10")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238_0\(81),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_4_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_0__G0_2_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2364_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_I_A2_3_RETO_0\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2473_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2470_RETO_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_10\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_14_10_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_10\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_51_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(51),
datain => N_80639,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_19_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(19),
datain => N_80671,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_0_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_11\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_15_10_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_11\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1_51_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(51),
datain => N_80639,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1_19_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(19),
datain => N_80671,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_1_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_12\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_16_10_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_12\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_2_51_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(51),
datain => N_80639,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_2_19_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(19),
datain => N_80671,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN39_ZERO_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000f33")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_5\(21),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_5\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_2_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_0\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_10\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_17_10_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_4\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_0\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_5_21_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_5\(21),
datain => N_80669,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_5_53_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_5\(53),
datain => N_80637,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN33_ZERO_0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f33ffffffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_6\(21),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_6\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_1_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_3_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_1\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_10\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_18_10_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_5\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_0\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_6_21_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_6\(21),
datain => N_80669,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_6_53_\: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_6\(53),
datain => N_80637,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_345_RNI9E6S: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"fefafefabafabafa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_644_RETO_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10927_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(49),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_27_S_0_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10918_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0_0\,
datag => N_55054_RETO_0);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_345: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10927_RETO_0\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10927\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_346: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(49),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(49),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_347: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_27_S_0_RETO_0\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_27_S_0\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_348: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10918_RETO_0\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10918\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_349: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(50),
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(50),
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_350: stratixii_lcell_ff port map (
regout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_RETO_0_0\,
datain => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_2748_0\,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_351: stratixii_lcell_ff port map (
regout => N_55054_RETO_0,
datain => N_55054,
clk => N_8,
	devpor => devpor,
	devclrn => devclrn,
	aclr => GND,
	aload => GND,
	sclr => GND,
	sload => GND,
	adatasdata => GND,
	ena => VCC);
GRLFPC2_0_COMB_V_STATE2_RNIP0GF: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff000f0000000000")
port map (
combout => \GRLFPC2_0.COMB.V.STATE0\,
dataf => \GRLFPC2_0.N_3422\,
datae => \GRLFPC2_0.N_1105\,
datad => \GRLFPC2_0.R.STATE\(1),
datac => \GRLFPC2_0.N_1213\);
GRLFPC2_0_COMB_UN1_MEXC_1_RNIBACJ1: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ecffefffa0a0a0a0")
port map (
combout => \GRLFPC2_0.N_1721\,
dataf => \GRLFPC2_0.COMB.V.STATE0\,
datae => \GRLFPC2_0.R.I.EXEC\,
datad => \GRLFPC2_0.R.I.V\,
datac => \GRLFPC2_0.V.I.EXEC_0_SQMUXA\,
datab => \GRLFPC2_0.N_1768\,
dataa => \GRLFPC2_0.N_1105\);
GRLFPC2_0_V_FSR_CEXC_0_SQMUXA0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"7f007f7f00000000")
port map (
combout => \GRLFPC2_0.V.FSR.CEXC_0_SQMUXA0\,
dataf => \GRLFPC2_0.R.I.V\,
datae => \GRLFPC2_0.R.X.LD\,
datad => \GRLFPC2_0.COMB.ISFPOP2_1\,
datac => N_395,
datab => N_396,
dataa => N_397);
GRLFPC2_0_V_FSR_AEXC_2_SQMUXA0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ff0000ffffffff")
port map (
combout => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA0\,
dataf => \GRLFPC2_0.R.I.V\,
datae => \GRLFPC2_0.R.X.LD\,
datad => \GRLFPC2_0.COMB.ISFPOP2_1\,
datac => \GRLFPC2_0.N_1132\);
GRLFPC2_0_V_FSR_AEXC_2_SQMUXA: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0303030300030303")
port map (
combout => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA\,
dataf => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA0\,
datae => \GRLFPC2_0.N_1720\,
datad => \GRLFPC2_0.N_1302\,
datac => \GRLFPC2_0.N_1517\,
datab => \GRLFPC2_0.N_1132\);
GRLFPC2_0_COMB_WREN125: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000002000000")
port map (
combout => \GRLFPC2_0.N_1586\,
dataf => \GRLFPC2_0.N_1721\,
datae => \GRLFPC2_0.N_1309\,
datad => \GRLFPC2_0.R.I.V\,
datac => \GRLFPC2_0.R.X.LD\,
datab => \GRLFPC2_0.COMB.ISFPOP2_1\,
dataa => \GRLFPC2_0.N_1720\);
GRLFPC2_0_V_FSR_CEXC_3_SQMUXA0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0fff0fffffffff")
port map (
combout => \GRLFPC2_0.V.FSR.CEXC_3_SQMUXA0\,
dataf => \GRLFPC2_0.N_1720\,
datae => \GRLFPC2_0.COMB.ISFPOP2_1\,
datad => \GRLFPC2_0.R.X.LD\,
datac => \GRLFPC2_0.R.I.V\);
GRLFPC2_0_V_FSR_CEXC_0_SQMUXA: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f0000000")
port map (
combout => \GRLFPC2_0.V.FSR.CEXC_0_SQMUXA\,
dataf => \GRLFPC2_0.N_1721\,
datae => \GRLFPC2_0.N_1309\,
datad => \GRLFPC2_0.N_1720\,
datac => \GRLFPC2_0.V.FSR.CEXC_0_SQMUXA0\);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV0_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"a0ff00c0a00000c0")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0\,
dataf => N_364,
datae => \GRLFPC2_0.V.FSR.CEXC_2_SQMUXA_0\,
datad => \GRLFPC2_0.N_1570\,
datac => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV_0\(1),
datab => \GRLFPC2_0.R.FSR.CEXC\(1),
dataa => \GRLFPC2_0.R.I.EXC\(1));
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV0_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"a0ff00c0a00000c0")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0_0\,
dataf => N_367,
datae => \GRLFPC2_0.V.FSR.CEXC_2_SQMUXA_0\,
datad => \GRLFPC2_0.N_1570\,
datac => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV_0\(4),
datab => \GRLFPC2_0.R.FSR.CEXC\(4),
dataa => \GRLFPC2_0.R.I.EXC\(4));
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV0_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"a0ff00c0a00000c0")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0_1\,
dataf => N_363,
datae => \GRLFPC2_0.V.FSR.CEXC_2_SQMUXA_0\,
datad => \GRLFPC2_0.N_1570\,
datac => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV_0\(0),
datab => \GRLFPC2_0.R.FSR.CEXC\(0),
dataa => \GRLFPC2_0.R.I.EXC\(0));
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV0_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"a0ff00c0a00000c0")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0_2\,
dataf => N_365,
datae => \GRLFPC2_0.V.FSR.CEXC_2_SQMUXA_0\,
datad => \GRLFPC2_0.N_1570\,
datac => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV_0\(2),
datab => \GRLFPC2_0.R.FSR.CEXC\(2),
dataa => \GRLFPC2_0.R.I.EXC\(2));
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV0_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"a0ff00c0a00000c0")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0_3\,
dataf => N_366,
datae => \GRLFPC2_0.V.FSR.CEXC_2_SQMUXA_0\,
datad => \GRLFPC2_0.N_1570\,
datac => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV_0\(3),
datab => \GRLFPC2_0.R.FSR.CEXC\(3),
dataa => \GRLFPC2_0.R.I.EXC\(3));
\GRLFPC2_0_V_FSR_FTT_1_IV_I_A3_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"e0a0e0a00000e0a0")
port map (
combout => \GRLFPC2_0.N_1570\,
dataf => \GRLFPC2_0.V.FSR.FTT_1_IV_I_A30\,
datae => \GRLFPC2_0.COMB.UN1_MEXC_1_0\,
datad => \GRLFPC2_0.R.I.EXEC\,
datac => \GRLFPC2_0.R.I.V\,
datab => \GRLFPC2_0.N_3422\,
dataa => \GRLFPC2_0.V.I.EXEC_0_SQMUXA\);
\GRLFPC2_0_V_FSR_FTT_1_IV_I_A30_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff8ff88f8f88888")
port map (
combout => \GRLFPC2_0.V.FSR.FTT_1_IV_I_A30\,
dataf => \GRLFPC2_0.R.I.EXC\(1),
datae => \GRLFPC2_0.R.I.EXC\(0),
datad => \GRLFPC2_0.R.FSR.TEM\(1),
datac => \GRLFPC2_0.R.FSR.TEM\(0),
datab => \GRLFPC2_0.R.FSR.TEM\(4),
dataa => \GRLFPC2_0.R.I.EXC\(4));
GRLFPC2_0_COMB_UN1_V_STATE0: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff000000ff")
port map (
combout => \GRLFPC2_0.COMB.UN1_V.STATE0\,
dataf => \GRLFPC2_0.N_1105\,
datae => \GRLFPC2_0.R.STATE\(0),
datad => \GRLFPC2_0.R.X.SEQERR\);
GRLFPC2_0_COMB_UN1_V_STATE: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"5555051500000000")
port map (
combout => \GRLFPC2_0.N_1302\,
dataf => \GRLFPC2_0.COMB.UN1_V.STATE0\,
datae => \GRLFPC2_0.N_1768\,
datad => \GRLFPC2_0.V.I.EXEC_0_SQMUXA\,
datac => \GRLFPC2_0.R.I.V\,
datab => \GRLFPC2_0.R.I.EXEC\,
dataa => \GRLFPC2_0.COMB.V.STATE0\);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV0_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0f0000ff0f")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV0\,
dataf => N_411,
datae => \GRLFPC2_0.N_1517\,
datad => N_371,
datac => \GRLFPC2_0.N_1132\);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV0_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0f0000ff0f")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV0_0\,
dataf => N_412,
datae => \GRLFPC2_0.N_1517\,
datad => N_372,
datac => \GRLFPC2_0.N_1132\);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV0_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0f0000ff0f")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV0_1\,
dataf => N_409,
datae => \GRLFPC2_0.N_1517\,
datad => N_369,
datac => \GRLFPC2_0.N_1132\);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV0_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0f0000ff0f")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV0_2\,
dataf => N_410,
datae => \GRLFPC2_0.N_1517\,
datad => N_370,
datac => \GRLFPC2_0.N_1132\);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV0_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0f0000ff0f")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV0_3\,
dataf => N_408,
datae => \GRLFPC2_0.N_1517\,
datad => N_368,
datac => \GRLFPC2_0.N_1132\);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV0_0_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000000000000")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV0_4\,
dataf => \GRLFPC2_0.V.FSR.CEXC_0_SQMUXA0\,
datae => \GRLFPC2_0.N_1720\,
datad => \GRLFPC2_0.N_1721\);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ddfcddaaddaaddaa")
port map (
combout => \GRLFPC2_0.R.FSR.AEXC_1_0_2__I0_I_0\,
dataf => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV0_4\,
datae => \GRLFPC2_0.N_1309\,
datad => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA\,
datac => \GRLFPC2_0.R.I.EXC\(2),
datab => \GRLFPC2_0.R.FSR.AEXC\(2),
dataa => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV0_2\);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV0_0_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000000000000")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV0_5\,
dataf => \GRLFPC2_0.V.FSR.CEXC_0_SQMUXA0\,
datae => \GRLFPC2_0.N_1720\,
datad => \GRLFPC2_0.N_1721\);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ddfcddaaddaaddaa")
port map (
combout => \GRLFPC2_0.R.FSR.AEXC_1_0_1__I0_I_1\,
dataf => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV0_5\,
datae => \GRLFPC2_0.N_1309\,
datad => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA\,
datac => \GRLFPC2_0.R.I.EXC\(1),
datab => \GRLFPC2_0.R.FSR.AEXC\(1),
dataa => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV0_1\);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV0_0_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000000000000")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV0_6\,
dataf => \GRLFPC2_0.V.FSR.CEXC_0_SQMUXA0\,
datae => \GRLFPC2_0.N_1720\,
datad => \GRLFPC2_0.N_1721\);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ddfcddaaddaaddaa")
port map (
combout => \GRLFPC2_0.R.FSR.AEXC_1_0_4__I0_I_0\,
dataf => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV0_6\,
datae => \GRLFPC2_0.N_1309\,
datad => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA\,
datac => \GRLFPC2_0.R.I.EXC\(4),
datab => \GRLFPC2_0.R.FSR.AEXC\(4),
dataa => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV0_0\);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV0_0_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000000000000")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV0_7\,
dataf => \GRLFPC2_0.V.FSR.CEXC_0_SQMUXA0\,
datae => \GRLFPC2_0.N_1720\,
datad => \GRLFPC2_0.N_1721\);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ddfcddaaddaaddaa")
port map (
combout => \GRLFPC2_0.R.FSR.AEXC_1_0_3__I0_I_1\,
dataf => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV0_7\,
datae => \GRLFPC2_0.N_1309\,
datad => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA\,
datac => \GRLFPC2_0.R.I.EXC\(3),
datab => \GRLFPC2_0.R.FSR.AEXC\(3),
dataa => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV0\);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV0_0_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff0000ff0000")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0_4\,
dataf => \GRLFPC2_0.N_1570\,
datae => \GRLFPC2_0.N_1309\,
datad => \GRLFPC2_0.V.FSR.CEXC_3_SQMUXA0\);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_3_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"eeeebbe2eeeebbaa")
port map (
combout => \GRLFPC2_0.R.FSR.CEXC_1_0_3__I0_I_0\,
dataf => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0_4\,
datae => \GRLFPC2_0.N_1517\,
datad => \GRLFPC2_0.N_1721\,
datac => \GRLFPC2_0.R.I.EXC\(3),
datab => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV_0\(3),
dataa => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0_3\);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV0_0_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000ff0000")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0_5\,
dataf => \GRLFPC2_0.N_1721\,
datae => \GRLFPC2_0.N_1309\,
datad => \GRLFPC2_0.V.FSR.CEXC_3_SQMUXA0\);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_2_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"eeeeeef3eeeeeebb")
port map (
combout => \GRLFPC2_0.R.FSR.CEXC_1_0_2__I0_I_1\,
dataf => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0_5\,
datae => \GRLFPC2_0.N_1570\,
datad => \GRLFPC2_0.N_1517\,
datac => \GRLFPC2_0.R.I.EXC\(2),
datab => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV_0\(2),
dataa => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0_2\);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV0_0_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000ff0000")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0_6\,
dataf => \GRLFPC2_0.N_1721\,
datae => \GRLFPC2_0.N_1309\,
datad => \GRLFPC2_0.V.FSR.CEXC_3_SQMUXA0\);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"eeeeeef3eeeeeebb")
port map (
combout => \GRLFPC2_0.R.FSR.CEXC_1_0_0__I0_I_1\,
dataf => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0_6\,
datae => \GRLFPC2_0.N_1570\,
datad => \GRLFPC2_0.N_1517\,
datac => \GRLFPC2_0.R.I.EXC\(0),
datab => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV_0\(0),
dataa => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0_1\);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_0_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffff0f0f0cccc")
port map (
combout => \GRLFPC2_0.R.FSR.AEXC_1_0_0__I0_I_0\,
dataf => \GRLFPC2_0.V.FSR.CEXC_0_SQMUXA\,
datae => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA\,
datad => \GRLFPC2_0.R.I.EXC\(0),
datac => \GRLFPC2_0.R.FSR.AEXC\(0),
datab => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV0_3\);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV0_0_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000ff0000")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0_7\,
dataf => \GRLFPC2_0.N_1721\,
datae => \GRLFPC2_0.N_1309\,
datad => \GRLFPC2_0.V.FSR.CEXC_3_SQMUXA0\);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_4_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"eeeeeef3eeeeeebb")
port map (
combout => \GRLFPC2_0.R.FSR.CEXC_1_0_4__I0_I_1\,
dataf => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0_7\,
datae => \GRLFPC2_0.N_1570\,
datad => \GRLFPC2_0.N_1517\,
datac => \GRLFPC2_0.R.I.EXC\(4),
datab => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV_0\(4),
dataa => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0_0\);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV0_0_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000ff0000")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0_8\,
dataf => \GRLFPC2_0.N_1721\,
datae => \GRLFPC2_0.N_1309\,
datad => \GRLFPC2_0.V.FSR.CEXC_3_SQMUXA0\);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_1_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"eeeeeef3eeeeeebb")
port map (
combout => \GRLFPC2_0.R.FSR.CEXC_1_0_1__I0_I_0\,
dataf => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0_8\,
datae => \GRLFPC2_0.N_1570\,
datad => \GRLFPC2_0.N_1517\,
datac => \GRLFPC2_0.R.I.EXC\(1),
datab => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV_0\(1),
dataa => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M20_108_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0aaf0f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M20\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
datad => \GRLFPC2_0.FPI.LDOP\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datab => \GRLFPC2_0.FPO.FRAC\(5),
dataa => \GRLFPC2_0.FPO.FRAC\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_108_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcfcfcfc0c0c0cfc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(108),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M20\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M20_110_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0aaf0f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M20_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
datad => \GRLFPC2_0.FPI.LDOP\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datab => \GRLFPC2_0.FPO.FRAC\(3),
dataa => \GRLFPC2_0.FPO.FRAC\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_110_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcfcfcfc0c0c0cfc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(110),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M20_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M20_111_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0aaf0f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M20_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
datad => \GRLFPC2_0.FPI.LDOP\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(2),
dataa => \GRLFPC2_0.FPO.FRAC\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_111_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcfcfcfc0c0c0cfc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(111),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M20_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M20_109_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0aaf0f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M20_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
datad => \GRLFPC2_0.FPI.LDOP\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datab => \GRLFPC2_0.FPO.FRAC\(4),
dataa => \GRLFPC2_0.FPO.FRAC\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_109_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcfcfcfc0c0c0cfc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(109),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M20_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M20_107_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0aaf0f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M20_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
datad => \GRLFPC2_0.FPI.LDOP\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
datab => \GRLFPC2_0.FPO.FRAC\(6),
dataa => \GRLFPC2_0.FPO.FRAC\(8));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_107_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcfcfcfc0c0c0cfc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(107),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M20_3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M20_102_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0aaf0f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M20_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
datad => \GRLFPC2_0.FPI.LDOP\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44),
datab => \GRLFPC2_0.FPO.FRAC\(11),
dataa => \GRLFPC2_0.FPO.FRAC\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_102_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcfcfcfc0c0c0cfc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(102),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M20_4\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M20_96_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0aaf0f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M20_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
datad => \GRLFPC2_0.FPI.LDOP\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
datab => \GRLFPC2_0.FPO.FRAC\(17),
dataa => \GRLFPC2_0.FPO.FRAC\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_96_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcfcfcfc0c0c0cfc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(96),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M20_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M20_93_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0aaf0f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M20_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
datad => \GRLFPC2_0.FPI.LDOP\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datab => \GRLFPC2_0.FPO.FRAC\(20),
dataa => \GRLFPC2_0.FPO.FRAC\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_93_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcfcfcfc0c0c0cfc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(93),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M20_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M20_112_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0aaf0f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M20_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
datad => \GRLFPC2_0.FPI.LDOP\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(1),
dataa => \GRLFPC2_0.FPO.FRAC\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_112_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcfcfcfc0c0c0cfc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(112),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M20_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_83_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffbefeb14100400")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(83),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M30\,
datae => \GRLFPC2_0.FPO.FRAC\(30),
datad => \GRLFPC2_0.FPO.FRAC\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_82_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffbefeb14100400")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(82),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M30_0\,
datae => \GRLFPC2_0.FPO.FRAC\(31),
datad => \GRLFPC2_0.FPO.FRAC\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M300_83_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cccaccaaccccaaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M300\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(4),
datad => \GRLFPC2_0.FPI.LDOP_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M30_83_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfffcffac0ffc0fa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M30\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M300\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4534_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M300_82_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cccaccaaccccaaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M300_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(4),
datad => \GRLFPC2_0.FPI.LDOP_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M30_82_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfffcffac0ffc0fa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M30_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M300_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4534_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_63_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffbefeb14100400")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(63),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M30_1\,
datae => \GRLFPC2_0.FPO.FRAC\(50),
datad => \GRLFPC2_0.FPO.FRAC\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_73_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffbefeb14100400")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(73),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M30_2\,
datae => \GRLFPC2_0.FPO.FRAC\(40),
datad => \GRLFPC2_0.FPO.FRAC\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_78_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffbefeb14100400")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(78),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M30_3\,
datae => \GRLFPC2_0.FPO.FRAC\(35),
datad => \GRLFPC2_0.FPO.FRAC\(37),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffbefeb14100400")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(61),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M30_4\,
datae => \GRLFPC2_0.FPO.FRAC\(52),
datad => \GRLFPC2_0.FPO.FRAC\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_69_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffbefeb14100400")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(69),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M30_5\,
datae => \GRLFPC2_0.FPO.FRAC\(44),
datad => \GRLFPC2_0.FPO.FRAC\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_75_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffbefeb14100400")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(75),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M30_6\,
datae => \GRLFPC2_0.FPO.FRAC\(38),
datad => \GRLFPC2_0.FPO.FRAC\(40),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_71_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffbefeb14100400")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(71),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M30_7\,
datae => \GRLFPC2_0.FPO.FRAC\(42),
datad => \GRLFPC2_0.FPO.FRAC\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M300_75_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"caaacaaacacaaaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M300_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(4),
datad => \GRLFPC2_0.FPI.LDOP_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4534_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M30_75_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfcfcacfc0c0cac0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M30_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M300_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(75),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M300_69_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"caaacaaacacaaaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M300_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(4),
datad => \GRLFPC2_0.FPI.LDOP_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4534_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M30_69_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfcfcacfc0c0cac0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M30_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M300_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(69),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M300_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"caaacaaacacaaaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M300_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(4),
datad => \GRLFPC2_0.FPI.LDOP_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4534_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M30_61_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfcfcacfc0c0cac0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M30_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M300_3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M300_78_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"caaacaaacacaaaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M300_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(4),
datad => \GRLFPC2_0.FPI.LDOP_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4534_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M30_78_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfcfcacfc0c0cac0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M30_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M300_4\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(78),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M300_73_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"caaacaaacacaaaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M300_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(4),
datad => \GRLFPC2_0.FPI.LDOP_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4534_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M30_73_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfcfcacfc0c0cac0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M30_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M300_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(73),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M300_63_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"caaacaaacacaaaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M300_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(4),
datad => \GRLFPC2_0.FPI.LDOP_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4534_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M30_63_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfcfcacfc0c0cac0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M30_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M300_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(63),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M300_71_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"caaacaaacacaaaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M300_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(4),
datad => \GRLFPC2_0.FPI.LDOP_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4534_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M30_71_\: stratixii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfcfcacfc0c0cac0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M30_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M300_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(71),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13));
N_7 <= RST_INTERNAL;
N_8 <= CLK_INTERNAL;
N_9 <= HOLDN_INTERNAL;
N_10 <= CPI_FLUSH_INTERNAL;
N_11 <= CPI_EXACK_INTERNAL;
N_12 <= CPI_A_RS1_INTERNAL;
N_13 <= CPI_A_RS1_INTERNAL_0;
N_14 <= CPI_A_RS1_INTERNAL_1;
N_16 <= CPI_A_RS1_INTERNAL_2;
N_17 <= CPI_A_RS1_INTERNAL_3;
N_18 <= CPI_D_PC_INTERNAL;
N_19 <= CPI_D_PC_INTERNAL_0;
N_20 <= CPI_D_PC_INTERNAL_1;
N_21 <= CPI_D_PC_INTERNAL_2;
N_22 <= CPI_D_PC_INTERNAL_3;
N_23 <= CPI_D_PC_INTERNAL_4;
N_24 <= CPI_D_PC_INTERNAL_5;
N_25 <= CPI_D_PC_INTERNAL_6;
N_26 <= CPI_D_PC_INTERNAL_7;
N_27 <= CPI_D_PC_INTERNAL_8;
N_28 <= CPI_D_PC_INTERNAL_9;
N_29 <= CPI_D_PC_INTERNAL_10;
N_30 <= CPI_D_PC_INTERNAL_11;
N_31 <= CPI_D_PC_INTERNAL_12;
N_32 <= CPI_D_PC_INTERNAL_13;
N_33 <= CPI_D_PC_INTERNAL_14;
N_34 <= CPI_D_PC_INTERNAL_15;
N_35 <= CPI_D_PC_INTERNAL_16;
N_36 <= CPI_D_PC_INTERNAL_17;
N_37 <= CPI_D_PC_INTERNAL_18;
N_38 <= CPI_D_PC_INTERNAL_19;
N_39 <= CPI_D_PC_INTERNAL_20;
N_40 <= CPI_D_PC_INTERNAL_21;
N_41 <= CPI_D_PC_INTERNAL_22;
N_42 <= CPI_D_PC_INTERNAL_23;
N_43 <= CPI_D_PC_INTERNAL_24;
N_44 <= CPI_D_PC_INTERNAL_25;
N_45 <= CPI_D_PC_INTERNAL_26;
N_46 <= CPI_D_PC_INTERNAL_27;
N_47 <= CPI_D_PC_INTERNAL_28;
N_48 <= CPI_D_PC_INTERNAL_29;
N_49 <= CPI_D_PC_INTERNAL_30;
N_50 <= CPI_D_INST_INTERNAL;
N_51 <= CPI_D_INST_INTERNAL_0;
N_52 <= CPI_D_INST_INTERNAL_1;
N_53 <= CPI_D_INST_INTERNAL_2;
N_54 <= CPI_D_INST_INTERNAL_3;
N_55 <= CPI_D_INST_INTERNAL_4;
N_56 <= CPI_D_INST_INTERNAL_5;
N_57 <= CPI_D_INST_INTERNAL_6;
N_58 <= CPI_D_INST_INTERNAL_7;
N_59 <= CPI_D_INST_INTERNAL_8;
N_60 <= CPI_D_INST_INTERNAL_9;
N_61 <= CPI_D_INST_INTERNAL_10;
N_62 <= CPI_D_INST_INTERNAL_11;
N_63 <= CPI_D_INST_INTERNAL_12;
N_64 <= CPI_D_INST_INTERNAL_13;
N_65 <= CPI_D_INST_INTERNAL_14;
N_66 <= CPI_D_INST_INTERNAL_15;
N_67 <= CPI_D_INST_INTERNAL_16;
N_68 <= CPI_D_INST_INTERNAL_17;
N_69 <= CPI_D_INST_INTERNAL_18;
N_70 <= CPI_D_INST_INTERNAL_19;
N_71 <= CPI_D_INST_INTERNAL_20;
N_72 <= CPI_D_INST_INTERNAL_21;
N_73 <= CPI_D_INST_INTERNAL_22;
N_74 <= CPI_D_INST_INTERNAL_23;
N_75 <= CPI_D_INST_INTERNAL_24;
N_76 <= CPI_D_INST_INTERNAL_25;
N_77 <= CPI_D_INST_INTERNAL_26;
N_78 <= CPI_D_INST_INTERNAL_27;
N_79 <= CPI_D_INST_INTERNAL_28;
N_80 <= CPI_D_INST_INTERNAL_29;
N_81 <= CPI_D_INST_INTERNAL_30;
N_82 <= CPI_D_CNT_INTERNAL;
N_83 <= CPI_D_CNT_INTERNAL_0;
N_84 <= CPI_D_TRAP_INTERNAL;
N_85 <= CPI_D_ANNUL_INTERNAL;
N_86 <= CPI_D_PV_INTERNAL;
N_87 <= CPI_A_PC_INTERNAL;
N_88 <= CPI_A_PC_INTERNAL_0;
N_89 <= CPI_A_PC_INTERNAL_1;
N_90 <= CPI_A_PC_INTERNAL_2;
N_91 <= CPI_A_PC_INTERNAL_3;
N_92 <= CPI_A_PC_INTERNAL_4;
N_93 <= CPI_A_PC_INTERNAL_5;
N_94 <= CPI_A_PC_INTERNAL_6;
N_95 <= CPI_A_PC_INTERNAL_7;
N_96 <= CPI_A_PC_INTERNAL_8;
N_97 <= CPI_A_PC_INTERNAL_9;
N_98 <= CPI_A_PC_INTERNAL_10;
N_99 <= CPI_A_PC_INTERNAL_11;
N_100 <= CPI_A_PC_INTERNAL_12;
N_101 <= CPI_A_PC_INTERNAL_13;
N_102 <= CPI_A_PC_INTERNAL_14;
N_103 <= CPI_A_PC_INTERNAL_15;
N_104 <= CPI_A_PC_INTERNAL_16;
N_105 <= CPI_A_PC_INTERNAL_17;
N_106 <= CPI_A_PC_INTERNAL_18;
N_107 <= CPI_A_PC_INTERNAL_19;
N_108 <= CPI_A_PC_INTERNAL_20;
N_109 <= CPI_A_PC_INTERNAL_21;
N_110 <= CPI_A_PC_INTERNAL_22;
N_111 <= CPI_A_PC_INTERNAL_23;
N_112 <= CPI_A_PC_INTERNAL_24;
N_113 <= CPI_A_PC_INTERNAL_25;
N_114 <= CPI_A_PC_INTERNAL_26;
N_115 <= CPI_A_PC_INTERNAL_27;
N_116 <= CPI_A_PC_INTERNAL_28;
N_117 <= CPI_A_PC_INTERNAL_29;
N_118 <= CPI_A_PC_INTERNAL_30;
N_119 <= CPI_A_INST_INTERNAL;
N_120 <= CPI_A_INST_INTERNAL_0;
N_121 <= CPI_A_INST_INTERNAL_1;
N_122 <= CPI_A_INST_INTERNAL_2;
N_123 <= CPI_A_INST_INTERNAL_3;
N_124 <= CPI_A_INST_INTERNAL_4;
N_125 <= CPI_A_INST_INTERNAL_5;
N_126 <= CPI_A_INST_INTERNAL_6;
N_127 <= CPI_A_INST_INTERNAL_7;
N_128 <= CPI_A_INST_INTERNAL_8;
N_129 <= CPI_A_INST_INTERNAL_9;
N_130 <= CPI_A_INST_INTERNAL_10;
N_131 <= CPI_A_INST_INTERNAL_11;
N_132 <= CPI_A_INST_INTERNAL_12;
N_133 <= CPI_A_INST_INTERNAL_13;
N_134 <= CPI_A_INST_INTERNAL_14;
N_135 <= CPI_A_INST_INTERNAL_15;
N_136 <= CPI_A_INST_INTERNAL_16;
N_137 <= CPI_A_INST_INTERNAL_17;
N_138 <= CPI_A_INST_INTERNAL_18;
N_139 <= CPI_A_INST_INTERNAL_19;
N_140 <= CPI_A_INST_INTERNAL_20;
N_141 <= CPI_A_INST_INTERNAL_21;
N_142 <= CPI_A_INST_INTERNAL_22;
N_143 <= CPI_A_INST_INTERNAL_23;
N_144 <= CPI_A_INST_INTERNAL_24;
N_145 <= CPI_A_INST_INTERNAL_25;
N_146 <= CPI_A_INST_INTERNAL_26;
N_147 <= CPI_A_INST_INTERNAL_27;
N_148 <= CPI_A_INST_INTERNAL_28;
N_149 <= CPI_A_INST_INTERNAL_29;
N_150 <= CPI_A_INST_INTERNAL_30;
N_151 <= CPI_A_CNT_INTERNAL;
N_152 <= CPI_A_CNT_INTERNAL_0;
N_153 <= CPI_A_TRAP_INTERNAL;
N_154 <= CPI_A_ANNUL_INTERNAL;
N_155 <= CPI_A_PV_INTERNAL;
N_156 <= CPI_E_PC_INTERNAL;
N_157 <= CPI_E_PC_INTERNAL_0;
N_158 <= CPI_E_PC_INTERNAL_1;
N_159 <= CPI_E_PC_INTERNAL_2;
N_160 <= CPI_E_PC_INTERNAL_3;
N_161 <= CPI_E_PC_INTERNAL_4;
N_162 <= CPI_E_PC_INTERNAL_5;
N_163 <= CPI_E_PC_INTERNAL_6;
N_164 <= CPI_E_PC_INTERNAL_7;
N_165 <= CPI_E_PC_INTERNAL_8;
N_166 <= CPI_E_PC_INTERNAL_9;
N_167 <= CPI_E_PC_INTERNAL_10;
N_168 <= CPI_E_PC_INTERNAL_11;
N_169 <= CPI_E_PC_INTERNAL_12;
N_170 <= CPI_E_PC_INTERNAL_13;
N_171 <= CPI_E_PC_INTERNAL_14;
N_172 <= CPI_E_PC_INTERNAL_15;
N_173 <= CPI_E_PC_INTERNAL_16;
N_174 <= CPI_E_PC_INTERNAL_17;
N_175 <= CPI_E_PC_INTERNAL_18;
N_176 <= CPI_E_PC_INTERNAL_19;
N_177 <= CPI_E_PC_INTERNAL_20;
N_178 <= CPI_E_PC_INTERNAL_21;
N_179 <= CPI_E_PC_INTERNAL_22;
N_180 <= CPI_E_PC_INTERNAL_23;
N_181 <= CPI_E_PC_INTERNAL_24;
N_182 <= CPI_E_PC_INTERNAL_25;
N_183 <= CPI_E_PC_INTERNAL_26;
N_184 <= CPI_E_PC_INTERNAL_27;
N_185 <= CPI_E_PC_INTERNAL_28;
N_186 <= CPI_E_PC_INTERNAL_29;
N_187 <= CPI_E_PC_INTERNAL_30;
N_188 <= CPI_E_INST_INTERNAL;
N_189 <= CPI_E_INST_INTERNAL_0;
N_190 <= CPI_E_INST_INTERNAL_1;
N_191 <= CPI_E_INST_INTERNAL_2;
N_192 <= CPI_E_INST_INTERNAL_3;
N_193 <= CPI_E_INST_INTERNAL_4;
N_194 <= CPI_E_INST_INTERNAL_5;
N_195 <= CPI_E_INST_INTERNAL_6;
N_196 <= CPI_E_INST_INTERNAL_7;
N_197 <= CPI_E_INST_INTERNAL_8;
N_198 <= CPI_E_INST_INTERNAL_9;
N_199 <= CPI_E_INST_INTERNAL_10;
N_200 <= CPI_E_INST_INTERNAL_11;
N_201 <= CPI_E_INST_INTERNAL_12;
N_202 <= CPI_E_INST_INTERNAL_13;
N_203 <= CPI_E_INST_INTERNAL_14;
N_204 <= CPI_E_INST_INTERNAL_15;
N_205 <= CPI_E_INST_INTERNAL_16;
N_206 <= CPI_E_INST_INTERNAL_17;
N_207 <= CPI_E_INST_INTERNAL_18;
N_208 <= CPI_E_INST_INTERNAL_19;
N_209 <= CPI_E_INST_INTERNAL_20;
N_210 <= CPI_E_INST_INTERNAL_21;
N_211 <= CPI_E_INST_INTERNAL_22;
N_212 <= CPI_E_INST_INTERNAL_23;
N_213 <= CPI_E_INST_INTERNAL_24;
N_214 <= CPI_E_INST_INTERNAL_25;
N_215 <= CPI_E_INST_INTERNAL_26;
N_216 <= CPI_E_INST_INTERNAL_27;
N_217 <= CPI_E_INST_INTERNAL_28;
N_218 <= CPI_E_INST_INTERNAL_29;
N_219 <= CPI_E_INST_INTERNAL_30;
N_220 <= CPI_E_CNT_INTERNAL;
N_221 <= CPI_E_CNT_INTERNAL_0;
N_222 <= CPI_E_TRAP_INTERNAL;
N_223 <= CPI_E_ANNUL_INTERNAL;
N_224 <= CPI_E_PV_INTERNAL;
N_225 <= CPI_M_PC_INTERNAL;
N_226 <= CPI_M_PC_INTERNAL_0;
N_227 <= CPI_M_PC_INTERNAL_1;
N_228 <= CPI_M_PC_INTERNAL_2;
N_229 <= CPI_M_PC_INTERNAL_3;
N_230 <= CPI_M_PC_INTERNAL_4;
N_231 <= CPI_M_PC_INTERNAL_5;
N_232 <= CPI_M_PC_INTERNAL_6;
N_233 <= CPI_M_PC_INTERNAL_7;
N_234 <= CPI_M_PC_INTERNAL_8;
N_235 <= CPI_M_PC_INTERNAL_9;
N_236 <= CPI_M_PC_INTERNAL_10;
N_237 <= CPI_M_PC_INTERNAL_11;
N_238 <= CPI_M_PC_INTERNAL_12;
N_239 <= CPI_M_PC_INTERNAL_13;
N_240 <= CPI_M_PC_INTERNAL_14;
N_241 <= CPI_M_PC_INTERNAL_15;
N_242 <= CPI_M_PC_INTERNAL_16;
N_243 <= CPI_M_PC_INTERNAL_17;
N_244 <= CPI_M_PC_INTERNAL_18;
N_245 <= CPI_M_PC_INTERNAL_19;
N_246 <= CPI_M_PC_INTERNAL_20;
N_247 <= CPI_M_PC_INTERNAL_21;
N_248 <= CPI_M_PC_INTERNAL_22;
N_249 <= CPI_M_PC_INTERNAL_23;
N_250 <= CPI_M_PC_INTERNAL_24;
N_251 <= CPI_M_PC_INTERNAL_25;
N_252 <= CPI_M_PC_INTERNAL_26;
N_253 <= CPI_M_PC_INTERNAL_27;
N_254 <= CPI_M_PC_INTERNAL_28;
N_255 <= CPI_M_PC_INTERNAL_29;
N_256 <= CPI_M_PC_INTERNAL_30;
N_257 <= CPI_M_INST_INTERNAL;
N_258 <= CPI_M_INST_INTERNAL_0;
N_259 <= CPI_M_INST_INTERNAL_1;
N_260 <= CPI_M_INST_INTERNAL_2;
N_261 <= CPI_M_INST_INTERNAL_3;
N_262 <= CPI_M_INST_INTERNAL_4;
N_263 <= CPI_M_INST_INTERNAL_5;
N_264 <= CPI_M_INST_INTERNAL_6;
N_265 <= CPI_M_INST_INTERNAL_7;
N_266 <= CPI_M_INST_INTERNAL_8;
N_267 <= CPI_M_INST_INTERNAL_9;
N_268 <= CPI_M_INST_INTERNAL_10;
N_269 <= CPI_M_INST_INTERNAL_11;
N_270 <= CPI_M_INST_INTERNAL_12;
N_271 <= CPI_M_INST_INTERNAL_13;
N_272 <= CPI_M_INST_INTERNAL_14;
N_273 <= CPI_M_INST_INTERNAL_15;
N_274 <= CPI_M_INST_INTERNAL_16;
N_275 <= CPI_M_INST_INTERNAL_17;
N_276 <= CPI_M_INST_INTERNAL_18;
N_277 <= CPI_M_INST_INTERNAL_19;
N_278 <= CPI_M_INST_INTERNAL_20;
N_279 <= CPI_M_INST_INTERNAL_21;
N_280 <= CPI_M_INST_INTERNAL_22;
N_281 <= CPI_M_INST_INTERNAL_23;
N_282 <= CPI_M_INST_INTERNAL_24;
N_283 <= CPI_M_INST_INTERNAL_25;
N_284 <= CPI_M_INST_INTERNAL_26;
N_285 <= CPI_M_INST_INTERNAL_27;
N_286 <= CPI_M_INST_INTERNAL_28;
N_287 <= CPI_M_INST_INTERNAL_29;
N_288 <= CPI_M_INST_INTERNAL_30;
N_289 <= CPI_M_CNT_INTERNAL;
N_290 <= CPI_M_CNT_INTERNAL_0;
N_291 <= CPI_M_TRAP_INTERNAL;
N_292 <= CPI_M_ANNUL_INTERNAL;
N_293 <= CPI_M_PV_INTERNAL;
N_294 <= CPI_X_PC_INTERNAL;
N_295 <= CPI_X_PC_INTERNAL_0;
N_296 <= CPI_X_PC_INTERNAL_1;
N_297 <= CPI_X_PC_INTERNAL_2;
N_298 <= CPI_X_PC_INTERNAL_3;
N_299 <= CPI_X_PC_INTERNAL_4;
N_300 <= CPI_X_PC_INTERNAL_5;
N_301 <= CPI_X_PC_INTERNAL_6;
N_302 <= CPI_X_PC_INTERNAL_7;
N_303 <= CPI_X_PC_INTERNAL_8;
N_304 <= CPI_X_PC_INTERNAL_9;
N_305 <= CPI_X_PC_INTERNAL_10;
N_306 <= CPI_X_PC_INTERNAL_11;
N_307 <= CPI_X_PC_INTERNAL_12;
N_308 <= CPI_X_PC_INTERNAL_13;
N_309 <= CPI_X_PC_INTERNAL_14;
N_310 <= CPI_X_PC_INTERNAL_15;
N_311 <= CPI_X_PC_INTERNAL_16;
N_312 <= CPI_X_PC_INTERNAL_17;
N_313 <= CPI_X_PC_INTERNAL_18;
N_314 <= CPI_X_PC_INTERNAL_19;
N_315 <= CPI_X_PC_INTERNAL_20;
N_316 <= CPI_X_PC_INTERNAL_21;
N_317 <= CPI_X_PC_INTERNAL_22;
N_318 <= CPI_X_PC_INTERNAL_23;
N_319 <= CPI_X_PC_INTERNAL_24;
N_320 <= CPI_X_PC_INTERNAL_25;
N_321 <= CPI_X_PC_INTERNAL_26;
N_322 <= CPI_X_PC_INTERNAL_27;
N_323 <= CPI_X_PC_INTERNAL_28;
N_324 <= CPI_X_PC_INTERNAL_29;
N_325 <= CPI_X_PC_INTERNAL_30;
N_326 <= CPI_X_INST_INTERNAL;
N_327 <= CPI_X_INST_INTERNAL_0;
N_328 <= CPI_X_INST_INTERNAL_1;
N_329 <= CPI_X_INST_INTERNAL_2;
N_330 <= CPI_X_INST_INTERNAL_3;
N_331 <= CPI_X_INST_INTERNAL_4;
N_332 <= CPI_X_INST_INTERNAL_5;
N_333 <= CPI_X_INST_INTERNAL_6;
N_334 <= CPI_X_INST_INTERNAL_7;
N_335 <= CPI_X_INST_INTERNAL_8;
N_336 <= CPI_X_INST_INTERNAL_9;
N_337 <= CPI_X_INST_INTERNAL_10;
N_338 <= CPI_X_INST_INTERNAL_11;
N_339 <= CPI_X_INST_INTERNAL_12;
N_340 <= CPI_X_INST_INTERNAL_13;
N_341 <= CPI_X_INST_INTERNAL_14;
N_342 <= CPI_X_INST_INTERNAL_15;
N_343 <= CPI_X_INST_INTERNAL_16;
N_344 <= CPI_X_INST_INTERNAL_17;
N_345 <= CPI_X_INST_INTERNAL_18;
N_346 <= CPI_X_INST_INTERNAL_19;
N_347 <= CPI_X_INST_INTERNAL_20;
N_348 <= CPI_X_INST_INTERNAL_21;
N_349 <= CPI_X_INST_INTERNAL_22;
N_350 <= CPI_X_INST_INTERNAL_23;
N_351 <= CPI_X_INST_INTERNAL_24;
N_352 <= CPI_X_INST_INTERNAL_25;
N_353 <= CPI_X_INST_INTERNAL_26;
N_354 <= CPI_X_INST_INTERNAL_27;
N_355 <= CPI_X_INST_INTERNAL_28;
N_356 <= CPI_X_INST_INTERNAL_29;
N_357 <= CPI_X_INST_INTERNAL_30;
N_358 <= CPI_X_CNT_INTERNAL;
N_359 <= CPI_X_CNT_INTERNAL_0;
N_360 <= CPI_X_TRAP_INTERNAL;
N_361 <= CPI_X_ANNUL_INTERNAL;
N_362 <= CPI_X_PV_INTERNAL;
N_363 <= CPI_LDDATA_INTERNAL;
N_364 <= CPI_LDDATA_INTERNAL_0;
N_365 <= CPI_LDDATA_INTERNAL_1;
N_366 <= CPI_LDDATA_INTERNAL_2;
N_367 <= CPI_LDDATA_INTERNAL_3;
N_368 <= CPI_LDDATA_INTERNAL_4;
N_369 <= CPI_LDDATA_INTERNAL_5;
N_370 <= CPI_LDDATA_INTERNAL_6;
N_371 <= CPI_LDDATA_INTERNAL_7;
N_372 <= CPI_LDDATA_INTERNAL_8;
N_373 <= CPI_LDDATA_INTERNAL_9;
N_374 <= CPI_LDDATA_INTERNAL_10;
N_375 <= CPI_LDDATA_INTERNAL_11;
N_376 <= CPI_LDDATA_INTERNAL_12;
N_377 <= CPI_LDDATA_INTERNAL_13;
N_378 <= CPI_LDDATA_INTERNAL_14;
N_379 <= CPI_LDDATA_INTERNAL_15;
N_380 <= CPI_LDDATA_INTERNAL_16;
N_381 <= CPI_LDDATA_INTERNAL_17;
N_382 <= CPI_LDDATA_INTERNAL_18;
N_383 <= CPI_LDDATA_INTERNAL_19;
N_384 <= CPI_LDDATA_INTERNAL_20;
N_385 <= CPI_LDDATA_INTERNAL_21;
N_386 <= CPI_LDDATA_INTERNAL_22;
N_387 <= CPI_LDDATA_INTERNAL_23;
N_388 <= CPI_LDDATA_INTERNAL_24;
N_389 <= CPI_LDDATA_INTERNAL_25;
N_390 <= CPI_LDDATA_INTERNAL_26;
N_391 <= CPI_LDDATA_INTERNAL_27;
N_392 <= CPI_LDDATA_INTERNAL_28;
N_393 <= CPI_LDDATA_INTERNAL_29;
N_394 <= CPI_LDDATA_INTERNAL_30;
N_395 <= CPI_DBG_ENABLE_INTERNAL;
N_396 <= CPI_DBG_WRITE_INTERNAL;
N_397 <= CPI_DBG_FSR_INTERNAL;
N_398 <= CPI_DBG_ADDR_INTERNAL;
N_399 <= CPI_DBG_ADDR_INTERNAL_0;
N_400 <= CPI_DBG_ADDR_INTERNAL_1;
N_401 <= CPI_DBG_ADDR_INTERNAL_2;
N_402 <= CPI_DBG_ADDR_INTERNAL_3;
N_403 <= CPI_DBG_DATA_INTERNAL;
N_404 <= CPI_DBG_DATA_INTERNAL_0;
N_405 <= CPI_DBG_DATA_INTERNAL_1;
N_406 <= CPI_DBG_DATA_INTERNAL_2;
N_407 <= CPI_DBG_DATA_INTERNAL_3;
N_408 <= CPI_DBG_DATA_INTERNAL_4;
N_409 <= CPI_DBG_DATA_INTERNAL_5;
N_410 <= CPI_DBG_DATA_INTERNAL_6;
N_411 <= CPI_DBG_DATA_INTERNAL_7;
N_412 <= CPI_DBG_DATA_INTERNAL_8;
N_413 <= CPI_DBG_DATA_INTERNAL_9;
N_414 <= CPI_DBG_DATA_INTERNAL_10;
N_415 <= CPI_DBG_DATA_INTERNAL_11;
N_416 <= CPI_DBG_DATA_INTERNAL_12;
N_417 <= CPI_DBG_DATA_INTERNAL_13;
N_418 <= CPI_DBG_DATA_INTERNAL_14;
N_419 <= CPI_DBG_DATA_INTERNAL_15;
N_420 <= CPI_DBG_DATA_INTERNAL_16;
N_421 <= CPI_DBG_DATA_INTERNAL_17;
N_422 <= CPI_DBG_DATA_INTERNAL_18;
N_423 <= CPI_DBG_DATA_INTERNAL_19;
N_424 <= CPI_DBG_DATA_INTERNAL_20;
N_425 <= CPI_DBG_DATA_INTERNAL_21;
N_426 <= CPI_DBG_DATA_INTERNAL_22;
N_427 <= CPI_DBG_DATA_INTERNAL_23;
N_428 <= CPI_DBG_DATA_INTERNAL_24;
N_429 <= CPI_DBG_DATA_INTERNAL_25;
N_430 <= CPI_DBG_DATA_INTERNAL_26;
N_431 <= CPI_DBG_DATA_INTERNAL_27;
N_432 <= CPI_DBG_DATA_INTERNAL_28;
N_433 <= CPI_DBG_DATA_INTERNAL_29;
N_434 <= CPI_DBG_DATA_INTERNAL_30;
N_0 <= CPO_DATAZ(0);
N_1_115 <= CPO_DATAZ(1);
N_2_116 <= CPO_DATAZ(2);
N_3_117 <= CPO_DATAZ(3);
N_4_118 <= CPO_DATAZ(4);
N_5_119 <= CPO_DATAZ(5);
N_6_120 <= CPO_DATAZ(6);
N_7_121 <= CPO_DATAZ(7);
N_8_122 <= CPO_DATAZ(8);
N_9_123 <= CPO_DATAZ(9);
N_10_124 <= CPO_DATAZ(10);
N_11_125 <= CPO_DATAZ(11);
N_12_126 <= CPO_DATAZ(12);
N_13_127 <= CPO_DATAZ(13);
N_14_128 <= CPO_DATAZ(14);
N_15_129 <= CPO_DATAZ(15);
N_16_130 <= CPO_DATAZ(16);
N_17_131 <= CPO_DATAZ(17);
N_18_132 <= CPO_DATAZ(18);
N_19_133 <= CPO_DATAZ(19);
N_20_134 <= CPO_DATAZ(20);
N_21_135 <= CPO_DATAZ(21);
N_22_136 <= CPO_DATAZ(22);
N_23_137 <= CPO_DATAZ(23);
N_24_138 <= CPO_DATAZ(24);
N_25_139 <= CPO_DATAZ(25);
N_26_140 <= CPO_DATAZ(26);
N_27_141 <= CPO_DATAZ(27);
N_28_142 <= CPO_DATAZ(28);
N_29_143 <= CPO_DATAZ(29);
N_30_144 <= CPO_DATAZ(30);
N_31_145 <= CPO_DATAZ(31);
N_32_146 <= CPO_EXCZ;
N_33_147 <= CPO_CCZ(0);
N_34_148 <= CPO_CCZ(1);
N_35_149 <= CPO_CCVZ;
N_36_150 <= CPO_LDLOCKZ;
N_37_151 <= CPO_HOLDNZ;
N_38_152 <= CPO_DBG_DATAZ(0);
N_39_153 <= CPO_DBG_DATAZ(1);
N_40_154 <= CPO_DBG_DATAZ(2);
N_41_155 <= CPO_DBG_DATAZ(3);
N_42_156 <= CPO_DBG_DATAZ(4);
N_43_157 <= CPO_DBG_DATAZ(5);
N_44_158 <= CPO_DBG_DATAZ(6);
N_45_159 <= CPO_DBG_DATAZ(7);
N_46_160 <= CPO_DBG_DATAZ(8);
N_47_161 <= CPO_DBG_DATAZ(9);
N_48_162 <= CPO_DBG_DATAZ(10);
N_49_163 <= CPO_DBG_DATAZ(11);
N_50_164 <= CPO_DBG_DATAZ(12);
N_51_165 <= CPO_DBG_DATAZ(13);
N_52_166 <= CPO_DBG_DATAZ(14);
N_53_167 <= CPO_DBG_DATAZ(15);
N_54_168 <= CPO_DBG_DATAZ(16);
N_55_169 <= CPO_DBG_DATAZ(17);
N_56_170 <= CPO_DBG_DATAZ(18);
N_57_171 <= CPO_DBG_DATAZ(19);
N_58_172 <= CPO_DBG_DATAZ(20);
N_59_173 <= CPO_DBG_DATAZ(21);
N_60_174 <= CPO_DBG_DATAZ(22);
N_61_175 <= CPO_DBG_DATAZ(23);
N_62_176 <= CPO_DBG_DATAZ(24);
N_63_177 <= CPO_DBG_DATAZ(25);
N_64_178 <= CPO_DBG_DATAZ(26);
N_65_179 <= CPO_DBG_DATAZ(27);
N_66_180 <= CPO_DBG_DATAZ(28);
N_67_181 <= CPO_DBG_DATAZ(29);
N_68_182 <= CPO_DBG_DATAZ(30);
N_69_183 <= CPO_DBG_DATAZ(31);
N_70_184 <= RFI2_RD1ADDRZ(0);
N_71_185 <= RFI2_RD1ADDRZ(1);
N_72_186 <= RFI2_RD1ADDRZ(2);
N_73_187 <= RFI2_RD1ADDRZ(3);
N_74_188 <= RFI2_RD2ADDRZ(0);
N_75_189 <= RFI2_RD2ADDRZ(1);
N_76_190 <= RFI2_RD2ADDRZ(2);
N_77_191 <= RFI2_RD2ADDRZ(3);
N_78_192 <= RFI2_WRADDRZ(0);
N_79_193 <= RFI2_WRADDRZ(1);
N_80_194 <= RFI2_WRADDRZ(2);
N_81_195 <= RFI2_WRADDRZ(3);
N_82_196 <= RFI1_WRDATAZ(0);
N_83_197 <= RFI1_WRDATAZ(1);
N_84_198 <= RFI1_WRDATAZ(2);
N_85_199 <= RFI1_WRDATAZ(3);
N_86_200 <= RFI1_WRDATAZ(4);
N_87_201 <= RFI1_WRDATAZ(5);
N_88_202 <= RFI1_WRDATAZ(6);
N_89_203 <= RFI1_WRDATAZ(7);
N_90_204 <= RFI1_WRDATAZ(8);
N_91_205 <= RFI1_WRDATAZ(9);
N_92_206 <= RFI1_WRDATAZ(10);
N_93_207 <= RFI1_WRDATAZ(11);
N_94_208 <= RFI1_WRDATAZ(12);
N_95_209 <= RFI1_WRDATAZ(13);
N_96_210 <= RFI1_WRDATAZ(14);
N_97_211 <= RFI1_WRDATAZ(15);
N_98_212 <= RFI1_WRDATAZ(16);
N_99_213 <= RFI1_WRDATAZ(17);
N_100_214 <= RFI1_WRDATAZ(18);
N_101_215 <= RFI1_WRDATAZ(19);
N_102_216 <= RFI1_WRDATAZ(20);
N_103_217 <= RFI1_WRDATAZ(21);
N_104_218 <= RFI1_WRDATAZ(22);
N_105_219 <= RFI1_WRDATAZ(23);
N_106_220 <= RFI1_WRDATAZ(24);
N_107_221 <= RFI1_WRDATAZ(25);
N_108_222 <= RFI1_WRDATAZ(26);
N_109_223 <= RFI1_WRDATAZ(27);
N_110_224 <= RFI1_WRDATAZ(28);
N_111_225 <= RFI1_WRDATAZ(29);
N_112_226 <= RFI1_WRDATAZ(30);
N_113_227 <= RFI1_WRDATAZ(31);
N_114_228 <= RFI1_REN1Z;
N_115_229 <= RFI1_REN2Z;
N_116_230 <= RFI1_WRENZ;
N_117_231 <= RFI2_RD1ADDRZ(0);
N_118_232 <= RFI2_RD1ADDRZ(1);
N_119_233 <= RFI2_RD1ADDRZ(2);
N_120_234 <= RFI2_RD1ADDRZ(3);
N_121_235 <= RFI2_RD2ADDRZ(0);
N_122_236 <= RFI2_RD2ADDRZ(1);
N_123_237 <= RFI2_RD2ADDRZ(2);
N_124_238 <= RFI2_RD2ADDRZ(3);
N_125_239 <= RFI2_WRADDRZ(0);
N_126_240 <= RFI2_WRADDRZ(1);
N_127_241 <= RFI2_WRADDRZ(2);
N_128_242 <= RFI2_WRADDRZ(3);
N_129_243 <= RFI2_WRDATAZ(0);
N_130_244 <= RFI2_WRDATAZ(1);
N_131_245 <= RFI2_WRDATAZ(2);
N_132_246 <= RFI2_WRDATAZ(3);
N_133_247 <= RFI2_WRDATAZ(4);
N_134_248 <= RFI2_WRDATAZ(5);
N_135_249 <= RFI2_WRDATAZ(6);
N_136_250 <= RFI2_WRDATAZ(7);
N_137_251 <= RFI2_WRDATAZ(8);
N_138_252 <= RFI2_WRDATAZ(9);
N_139_253 <= RFI2_WRDATAZ(10);
N_140_254 <= RFI2_WRDATAZ(11);
N_141_255 <= RFI2_WRDATAZ(12);
N_142_256 <= RFI2_WRDATAZ(13);
N_143_257 <= RFI2_WRDATAZ(14);
N_144_258 <= RFI2_WRDATAZ(15);
N_145_259 <= RFI2_WRDATAZ(16);
N_146_260 <= RFI2_WRDATAZ(17);
N_147_261 <= RFI2_WRDATAZ(18);
N_148_262 <= RFI2_WRDATAZ(19);
N_149_263 <= RFI2_WRDATAZ(20);
N_150_264 <= RFI2_WRDATAZ(21);
N_151_265 <= RFI2_WRDATAZ(22);
N_152_266 <= RFI2_WRDATAZ(23);
N_153_267 <= RFI2_WRDATAZ(24);
N_154_268 <= RFI2_WRDATAZ(25);
N_155_269 <= RFI2_WRDATAZ(26);
N_156_270 <= RFI2_WRDATAZ(27);
N_157_271 <= RFI2_WRDATAZ(28);
N_158_272 <= RFI2_WRDATAZ(29);
N_159_273 <= RFI2_WRDATAZ(30);
N_160_274 <= RFI2_WRDATAZ(31);
N_161_275 <= RFI2_REN1Z;
N_162_276 <= RFI2_REN2Z;
N_163_277 <= RFI2_WRENZ;
N_599 <= RFO1_DATA1_INTERNAL;
N_600 <= RFO1_DATA1_INTERNAL_0;
N_601 <= RFO1_DATA1_INTERNAL_1;
N_602 <= RFO1_DATA1_INTERNAL_2;
N_603 <= RFO1_DATA1_INTERNAL_3;
N_604 <= RFO1_DATA1_INTERNAL_4;
N_605 <= RFO1_DATA1_INTERNAL_5;
N_606 <= RFO1_DATA1_INTERNAL_6;
N_607 <= RFO1_DATA1_INTERNAL_7;
N_608 <= RFO1_DATA1_INTERNAL_8;
N_609 <= RFO1_DATA1_INTERNAL_9;
N_610 <= RFO1_DATA1_INTERNAL_10;
N_611 <= RFO1_DATA1_INTERNAL_11;
N_612 <= RFO1_DATA1_INTERNAL_12;
N_613 <= RFO1_DATA1_INTERNAL_13;
N_614 <= RFO1_DATA1_INTERNAL_14;
N_615 <= RFO1_DATA1_INTERNAL_15;
N_616 <= RFO1_DATA1_INTERNAL_16;
N_617 <= RFO1_DATA1_INTERNAL_17;
N_618 <= RFO1_DATA1_INTERNAL_18;
N_619 <= RFO1_DATA1_INTERNAL_19;
N_620 <= RFO1_DATA1_INTERNAL_20;
N_621 <= RFO1_DATA1_INTERNAL_21;
N_622 <= RFO1_DATA1_INTERNAL_22;
N_623 <= RFO1_DATA1_INTERNAL_23;
N_624 <= RFO1_DATA1_INTERNAL_24;
N_625 <= RFO1_DATA1_INTERNAL_25;
N_626 <= RFO1_DATA1_INTERNAL_26;
N_627 <= RFO1_DATA1_INTERNAL_27;
N_628 <= RFO1_DATA1_INTERNAL_28;
N_629 <= RFO1_DATA1_INTERNAL_29;
N_630 <= RFO1_DATA1_INTERNAL_30;
N_631 <= RFO1_DATA2_INTERNAL;
N_632 <= RFO1_DATA2_INTERNAL_0;
N_633 <= RFO1_DATA2_INTERNAL_1;
N_634 <= RFO1_DATA2_INTERNAL_2;
N_635 <= RFO1_DATA2_INTERNAL_3;
N_636 <= RFO1_DATA2_INTERNAL_4;
N_637 <= RFO1_DATA2_INTERNAL_5;
N_638 <= RFO1_DATA2_INTERNAL_6;
N_639 <= RFO1_DATA2_INTERNAL_7;
N_640 <= RFO1_DATA2_INTERNAL_8;
N_641 <= RFO1_DATA2_INTERNAL_9;
N_642 <= RFO1_DATA2_INTERNAL_10;
N_643 <= RFO1_DATA2_INTERNAL_11;
N_644 <= RFO1_DATA2_INTERNAL_12;
N_645 <= RFO1_DATA2_INTERNAL_13;
N_646 <= RFO1_DATA2_INTERNAL_14;
N_647 <= RFO1_DATA2_INTERNAL_15;
N_648 <= RFO1_DATA2_INTERNAL_16;
N_649 <= RFO1_DATA2_INTERNAL_17;
N_650 <= RFO1_DATA2_INTERNAL_18;
N_651 <= RFO1_DATA2_INTERNAL_19;
N_652 <= RFO1_DATA2_INTERNAL_20;
N_653 <= RFO1_DATA2_INTERNAL_21;
N_654 <= RFO1_DATA2_INTERNAL_22;
N_655 <= RFO1_DATA2_INTERNAL_23;
N_656 <= RFO1_DATA2_INTERNAL_24;
N_657 <= RFO1_DATA2_INTERNAL_25;
N_658 <= RFO1_DATA2_INTERNAL_26;
N_659 <= RFO1_DATA2_INTERNAL_27;
N_660 <= RFO1_DATA2_INTERNAL_28;
N_661 <= RFO1_DATA2_INTERNAL_29;
N_662 <= RFO1_DATA2_INTERNAL_30;
N_663 <= RFO2_DATA1_INTERNAL;
N_664 <= RFO2_DATA1_INTERNAL_0;
N_665 <= RFO2_DATA1_INTERNAL_1;
N_666 <= RFO2_DATA1_INTERNAL_2;
N_667 <= RFO2_DATA1_INTERNAL_3;
N_668 <= RFO2_DATA1_INTERNAL_4;
N_669 <= RFO2_DATA1_INTERNAL_5;
N_670 <= RFO2_DATA1_INTERNAL_6;
N_671 <= RFO2_DATA1_INTERNAL_7;
N_672 <= RFO2_DATA1_INTERNAL_8;
N_673 <= RFO2_DATA1_INTERNAL_9;
N_674 <= RFO2_DATA1_INTERNAL_10;
N_675 <= RFO2_DATA1_INTERNAL_11;
N_676 <= RFO2_DATA1_INTERNAL_12;
N_677 <= RFO2_DATA1_INTERNAL_13;
N_678 <= RFO2_DATA1_INTERNAL_14;
N_679 <= RFO2_DATA1_INTERNAL_15;
N_680 <= RFO2_DATA1_INTERNAL_16;
N_681 <= RFO2_DATA1_INTERNAL_17;
N_682 <= RFO2_DATA1_INTERNAL_18;
N_683 <= RFO2_DATA1_INTERNAL_19;
N_684 <= RFO2_DATA1_INTERNAL_20;
N_685 <= RFO2_DATA1_INTERNAL_21;
N_686 <= RFO2_DATA1_INTERNAL_22;
N_687 <= RFO2_DATA1_INTERNAL_23;
N_688 <= RFO2_DATA1_INTERNAL_24;
N_689 <= RFO2_DATA1_INTERNAL_25;
N_690 <= RFO2_DATA1_INTERNAL_26;
N_691 <= RFO2_DATA1_INTERNAL_27;
N_692 <= RFO2_DATA1_INTERNAL_28;
N_693 <= RFO2_DATA1_INTERNAL_29;
N_694 <= RFO2_DATA1_INTERNAL_30;
N_695 <= RFO2_DATA2_INTERNAL;
N_696 <= RFO2_DATA2_INTERNAL_0;
N_697 <= RFO2_DATA2_INTERNAL_1;
N_698 <= RFO2_DATA2_INTERNAL_2;
N_699 <= RFO2_DATA2_INTERNAL_3;
N_700 <= RFO2_DATA2_INTERNAL_4;
N_701 <= RFO2_DATA2_INTERNAL_5;
N_702 <= RFO2_DATA2_INTERNAL_6;
N_703 <= RFO2_DATA2_INTERNAL_7;
N_704 <= RFO2_DATA2_INTERNAL_8;
N_705 <= RFO2_DATA2_INTERNAL_9;
N_706 <= RFO2_DATA2_INTERNAL_10;
N_707 <= RFO2_DATA2_INTERNAL_11;
N_708 <= RFO2_DATA2_INTERNAL_12;
N_709 <= RFO2_DATA2_INTERNAL_13;
N_710 <= RFO2_DATA2_INTERNAL_14;
N_711 <= RFO2_DATA2_INTERNAL_15;
N_712 <= RFO2_DATA2_INTERNAL_16;
N_713 <= RFO2_DATA2_INTERNAL_17;
N_714 <= RFO2_DATA2_INTERNAL_18;
N_715 <= RFO2_DATA2_INTERNAL_19;
N_716 <= RFO2_DATA2_INTERNAL_20;
N_717 <= RFO2_DATA2_INTERNAL_21;
N_718 <= RFO2_DATA2_INTERNAL_22;
N_719 <= RFO2_DATA2_INTERNAL_23;
N_720 <= RFO2_DATA2_INTERNAL_24;
N_721 <= RFO2_DATA2_INTERNAL_25;
N_722 <= RFO2_DATA2_INTERNAL_26;
N_723 <= RFO2_DATA2_INTERNAL_27;
N_724 <= RFO2_DATA2_INTERNAL_28;
N_725 <= RFO2_DATA2_INTERNAL_29;
N_726 <= RFO2_DATA2_INTERNAL_30;
cpo_data(0) <= N_0;
cpo_data(1) <= N_1_115;
cpo_data(2) <= N_2_116;
cpo_data(3) <= N_3_117;
cpo_data(4) <= N_4_118;
cpo_data(5) <= N_5_119;
cpo_data(6) <= N_6_120;
cpo_data(7) <= N_7_121;
cpo_data(8) <= N_8_122;
cpo_data(9) <= N_9_123;
cpo_data(10) <= N_10_124;
cpo_data(11) <= N_11_125;
cpo_data(12) <= N_12_126;
cpo_data(13) <= N_13_127;
cpo_data(14) <= N_14_128;
cpo_data(15) <= N_15_129;
cpo_data(16) <= N_16_130;
cpo_data(17) <= N_17_131;
cpo_data(18) <= N_18_132;
cpo_data(19) <= N_19_133;
cpo_data(20) <= N_20_134;
cpo_data(21) <= N_21_135;
cpo_data(22) <= N_22_136;
cpo_data(23) <= N_23_137;
cpo_data(24) <= N_24_138;
cpo_data(25) <= N_25_139;
cpo_data(26) <= N_26_140;
cpo_data(27) <= N_27_141;
cpo_data(28) <= N_28_142;
cpo_data(29) <= N_29_143;
cpo_data(30) <= N_30_144;
cpo_data(31) <= N_31_145;
cpo_exc <= N_32_146;
cpo_cc(0) <= N_33_147;
cpo_cc(1) <= N_34_148;
cpo_ccv <= N_35_149;
cpo_ldlock <= N_36_150;
cpo_holdn <= N_37_151;
cpo_dbg_data(0) <= N_38_152;
cpo_dbg_data(1) <= N_39_153;
cpo_dbg_data(2) <= N_40_154;
cpo_dbg_data(3) <= N_41_155;
cpo_dbg_data(4) <= N_42_156;
cpo_dbg_data(5) <= N_43_157;
cpo_dbg_data(6) <= N_44_158;
cpo_dbg_data(7) <= N_45_159;
cpo_dbg_data(8) <= N_46_160;
cpo_dbg_data(9) <= N_47_161;
cpo_dbg_data(10) <= N_48_162;
cpo_dbg_data(11) <= N_49_163;
cpo_dbg_data(12) <= N_50_164;
cpo_dbg_data(13) <= N_51_165;
cpo_dbg_data(14) <= N_52_166;
cpo_dbg_data(15) <= N_53_167;
cpo_dbg_data(16) <= N_54_168;
cpo_dbg_data(17) <= N_55_169;
cpo_dbg_data(18) <= N_56_170;
cpo_dbg_data(19) <= N_57_171;
cpo_dbg_data(20) <= N_58_172;
cpo_dbg_data(21) <= N_59_173;
cpo_dbg_data(22) <= N_60_174;
cpo_dbg_data(23) <= N_61_175;
cpo_dbg_data(24) <= N_62_176;
cpo_dbg_data(25) <= N_63_177;
cpo_dbg_data(26) <= N_64_178;
cpo_dbg_data(27) <= N_65_179;
cpo_dbg_data(28) <= N_66_180;
cpo_dbg_data(29) <= N_67_181;
cpo_dbg_data(30) <= N_68_182;
cpo_dbg_data(31) <= N_69_183;
rfi1_rd1addr(0) <= N_70_184;
rfi1_rd1addr(1) <= N_71_185;
rfi1_rd1addr(2) <= N_72_186;
rfi1_rd1addr(3) <= N_73_187;
rfi1_rd2addr(0) <= N_74_188;
rfi1_rd2addr(1) <= N_75_189;
rfi1_rd2addr(2) <= N_76_190;
rfi1_rd2addr(3) <= N_77_191;
rfi1_wraddr(0) <= N_78_192;
rfi1_wraddr(1) <= N_79_193;
rfi1_wraddr(2) <= N_80_194;
rfi1_wraddr(3) <= N_81_195;
rfi1_wrdata(0) <= N_82_196;
rfi1_wrdata(1) <= N_83_197;
rfi1_wrdata(2) <= N_84_198;
rfi1_wrdata(3) <= N_85_199;
rfi1_wrdata(4) <= N_86_200;
rfi1_wrdata(5) <= N_87_201;
rfi1_wrdata(6) <= N_88_202;
rfi1_wrdata(7) <= N_89_203;
rfi1_wrdata(8) <= N_90_204;
rfi1_wrdata(9) <= N_91_205;
rfi1_wrdata(10) <= N_92_206;
rfi1_wrdata(11) <= N_93_207;
rfi1_wrdata(12) <= N_94_208;
rfi1_wrdata(13) <= N_95_209;
rfi1_wrdata(14) <= N_96_210;
rfi1_wrdata(15) <= N_97_211;
rfi1_wrdata(16) <= N_98_212;
rfi1_wrdata(17) <= N_99_213;
rfi1_wrdata(18) <= N_100_214;
rfi1_wrdata(19) <= N_101_215;
rfi1_wrdata(20) <= N_102_216;
rfi1_wrdata(21) <= N_103_217;
rfi1_wrdata(22) <= N_104_218;
rfi1_wrdata(23) <= N_105_219;
rfi1_wrdata(24) <= N_106_220;
rfi1_wrdata(25) <= N_107_221;
rfi1_wrdata(26) <= N_108_222;
rfi1_wrdata(27) <= N_109_223;
rfi1_wrdata(28) <= N_110_224;
rfi1_wrdata(29) <= N_111_225;
rfi1_wrdata(30) <= N_112_226;
rfi1_wrdata(31) <= N_113_227;
rfi1_ren1 <= N_114_228;
rfi1_ren2 <= N_115_229;
rfi1_wren <= N_116_230;
rfi2_rd1addr(0) <= N_117_231;
rfi2_rd1addr(1) <= N_118_232;
rfi2_rd1addr(2) <= N_119_233;
rfi2_rd1addr(3) <= N_120_234;
rfi2_rd2addr(0) <= N_121_235;
rfi2_rd2addr(1) <= N_122_236;
rfi2_rd2addr(2) <= N_123_237;
rfi2_rd2addr(3) <= N_124_238;
rfi2_wraddr(0) <= N_125_239;
rfi2_wraddr(1) <= N_126_240;
rfi2_wraddr(2) <= N_127_241;
rfi2_wraddr(3) <= N_128_242;
rfi2_wrdata(0) <= N_129_243;
rfi2_wrdata(1) <= N_130_244;
rfi2_wrdata(2) <= N_131_245;
rfi2_wrdata(3) <= N_132_246;
rfi2_wrdata(4) <= N_133_247;
rfi2_wrdata(5) <= N_134_248;
rfi2_wrdata(6) <= N_135_249;
rfi2_wrdata(7) <= N_136_250;
rfi2_wrdata(8) <= N_137_251;
rfi2_wrdata(9) <= N_138_252;
rfi2_wrdata(10) <= N_139_253;
rfi2_wrdata(11) <= N_140_254;
rfi2_wrdata(12) <= N_141_255;
rfi2_wrdata(13) <= N_142_256;
rfi2_wrdata(14) <= N_143_257;
rfi2_wrdata(15) <= N_144_258;
rfi2_wrdata(16) <= N_145_259;
rfi2_wrdata(17) <= N_146_260;
rfi2_wrdata(18) <= N_147_261;
rfi2_wrdata(19) <= N_148_262;
rfi2_wrdata(20) <= N_149_263;
rfi2_wrdata(21) <= N_150_264;
rfi2_wrdata(22) <= N_151_265;
rfi2_wrdata(23) <= N_152_266;
rfi2_wrdata(24) <= N_153_267;
rfi2_wrdata(25) <= N_154_268;
rfi2_wrdata(26) <= N_155_269;
rfi2_wrdata(27) <= N_156_270;
rfi2_wrdata(28) <= N_157_271;
rfi2_wrdata(29) <= N_158_272;
rfi2_wrdata(30) <= N_159_273;
rfi2_wrdata(31) <= N_160_274;
rfi2_ren1 <= N_161_275;
rfi2_ren2 <= N_162_276;
rfi2_wren <= N_163_277;
RST_INTERNAL <= rst;
CLK_INTERNAL <= clk;
HOLDN_INTERNAL <= holdn;
CPI_FLUSH_INTERNAL <= cpi_flush;
CPI_EXACK_INTERNAL <= cpi_exack;
CPI_A_RS1_INTERNAL <= cpi_a_rs1(0);
CPI_A_RS1_INTERNAL_0 <= cpi_a_rs1(1);
CPI_A_RS1_INTERNAL_1 <= cpi_a_rs1(2);
CPI_A_RS1_INTERNAL_2 <= cpi_a_rs1(3);
CPI_A_RS1_INTERNAL_3 <= cpi_a_rs1(4);
CPI_D_PC_INTERNAL <= cpi_d_pc(0);
CPI_D_PC_INTERNAL_0 <= cpi_d_pc(1);
CPI_D_PC_INTERNAL_1 <= cpi_d_pc(2);
CPI_D_PC_INTERNAL_2 <= cpi_d_pc(3);
CPI_D_PC_INTERNAL_3 <= cpi_d_pc(4);
CPI_D_PC_INTERNAL_4 <= cpi_d_pc(5);
CPI_D_PC_INTERNAL_5 <= cpi_d_pc(6);
CPI_D_PC_INTERNAL_6 <= cpi_d_pc(7);
CPI_D_PC_INTERNAL_7 <= cpi_d_pc(8);
CPI_D_PC_INTERNAL_8 <= cpi_d_pc(9);
CPI_D_PC_INTERNAL_9 <= cpi_d_pc(10);
CPI_D_PC_INTERNAL_10 <= cpi_d_pc(11);
CPI_D_PC_INTERNAL_11 <= cpi_d_pc(12);
CPI_D_PC_INTERNAL_12 <= cpi_d_pc(13);
CPI_D_PC_INTERNAL_13 <= cpi_d_pc(14);
CPI_D_PC_INTERNAL_14 <= cpi_d_pc(15);
CPI_D_PC_INTERNAL_15 <= cpi_d_pc(16);
CPI_D_PC_INTERNAL_16 <= cpi_d_pc(17);
CPI_D_PC_INTERNAL_17 <= cpi_d_pc(18);
CPI_D_PC_INTERNAL_18 <= cpi_d_pc(19);
CPI_D_PC_INTERNAL_19 <= cpi_d_pc(20);
CPI_D_PC_INTERNAL_20 <= cpi_d_pc(21);
CPI_D_PC_INTERNAL_21 <= cpi_d_pc(22);
CPI_D_PC_INTERNAL_22 <= cpi_d_pc(23);
CPI_D_PC_INTERNAL_23 <= cpi_d_pc(24);
CPI_D_PC_INTERNAL_24 <= cpi_d_pc(25);
CPI_D_PC_INTERNAL_25 <= cpi_d_pc(26);
CPI_D_PC_INTERNAL_26 <= cpi_d_pc(27);
CPI_D_PC_INTERNAL_27 <= cpi_d_pc(28);
CPI_D_PC_INTERNAL_28 <= cpi_d_pc(29);
CPI_D_PC_INTERNAL_29 <= cpi_d_pc(30);
CPI_D_PC_INTERNAL_30 <= cpi_d_pc(31);
CPI_D_INST_INTERNAL <= cpi_d_inst(0);
CPI_D_INST_INTERNAL_0 <= cpi_d_inst(1);
CPI_D_INST_INTERNAL_1 <= cpi_d_inst(2);
CPI_D_INST_INTERNAL_2 <= cpi_d_inst(3);
CPI_D_INST_INTERNAL_3 <= cpi_d_inst(4);
CPI_D_INST_INTERNAL_4 <= cpi_d_inst(5);
CPI_D_INST_INTERNAL_5 <= cpi_d_inst(6);
CPI_D_INST_INTERNAL_6 <= cpi_d_inst(7);
CPI_D_INST_INTERNAL_7 <= cpi_d_inst(8);
CPI_D_INST_INTERNAL_8 <= cpi_d_inst(9);
CPI_D_INST_INTERNAL_9 <= cpi_d_inst(10);
CPI_D_INST_INTERNAL_10 <= cpi_d_inst(11);
CPI_D_INST_INTERNAL_11 <= cpi_d_inst(12);
CPI_D_INST_INTERNAL_12 <= cpi_d_inst(13);
CPI_D_INST_INTERNAL_13 <= cpi_d_inst(14);
CPI_D_INST_INTERNAL_14 <= cpi_d_inst(15);
CPI_D_INST_INTERNAL_15 <= cpi_d_inst(16);
CPI_D_INST_INTERNAL_16 <= cpi_d_inst(17);
CPI_D_INST_INTERNAL_17 <= cpi_d_inst(18);
CPI_D_INST_INTERNAL_18 <= cpi_d_inst(19);
CPI_D_INST_INTERNAL_19 <= cpi_d_inst(20);
CPI_D_INST_INTERNAL_20 <= cpi_d_inst(21);
CPI_D_INST_INTERNAL_21 <= cpi_d_inst(22);
CPI_D_INST_INTERNAL_22 <= cpi_d_inst(23);
CPI_D_INST_INTERNAL_23 <= cpi_d_inst(24);
CPI_D_INST_INTERNAL_24 <= cpi_d_inst(25);
CPI_D_INST_INTERNAL_25 <= cpi_d_inst(26);
CPI_D_INST_INTERNAL_26 <= cpi_d_inst(27);
CPI_D_INST_INTERNAL_27 <= cpi_d_inst(28);
CPI_D_INST_INTERNAL_28 <= cpi_d_inst(29);
CPI_D_INST_INTERNAL_29 <= cpi_d_inst(30);
CPI_D_INST_INTERNAL_30 <= cpi_d_inst(31);
CPI_D_CNT_INTERNAL <= cpi_d_cnt(0);
CPI_D_CNT_INTERNAL_0 <= cpi_d_cnt(1);
CPI_D_TRAP_INTERNAL <= cpi_d_trap;
CPI_D_ANNUL_INTERNAL <= cpi_d_annul;
CPI_D_PV_INTERNAL <= cpi_d_pv;
CPI_A_PC_INTERNAL <= cpi_a_pc(0);
CPI_A_PC_INTERNAL_0 <= cpi_a_pc(1);
CPI_A_PC_INTERNAL_1 <= cpi_a_pc(2);
CPI_A_PC_INTERNAL_2 <= cpi_a_pc(3);
CPI_A_PC_INTERNAL_3 <= cpi_a_pc(4);
CPI_A_PC_INTERNAL_4 <= cpi_a_pc(5);
CPI_A_PC_INTERNAL_5 <= cpi_a_pc(6);
CPI_A_PC_INTERNAL_6 <= cpi_a_pc(7);
CPI_A_PC_INTERNAL_7 <= cpi_a_pc(8);
CPI_A_PC_INTERNAL_8 <= cpi_a_pc(9);
CPI_A_PC_INTERNAL_9 <= cpi_a_pc(10);
CPI_A_PC_INTERNAL_10 <= cpi_a_pc(11);
CPI_A_PC_INTERNAL_11 <= cpi_a_pc(12);
CPI_A_PC_INTERNAL_12 <= cpi_a_pc(13);
CPI_A_PC_INTERNAL_13 <= cpi_a_pc(14);
CPI_A_PC_INTERNAL_14 <= cpi_a_pc(15);
CPI_A_PC_INTERNAL_15 <= cpi_a_pc(16);
CPI_A_PC_INTERNAL_16 <= cpi_a_pc(17);
CPI_A_PC_INTERNAL_17 <= cpi_a_pc(18);
CPI_A_PC_INTERNAL_18 <= cpi_a_pc(19);
CPI_A_PC_INTERNAL_19 <= cpi_a_pc(20);
CPI_A_PC_INTERNAL_20 <= cpi_a_pc(21);
CPI_A_PC_INTERNAL_21 <= cpi_a_pc(22);
CPI_A_PC_INTERNAL_22 <= cpi_a_pc(23);
CPI_A_PC_INTERNAL_23 <= cpi_a_pc(24);
CPI_A_PC_INTERNAL_24 <= cpi_a_pc(25);
CPI_A_PC_INTERNAL_25 <= cpi_a_pc(26);
CPI_A_PC_INTERNAL_26 <= cpi_a_pc(27);
CPI_A_PC_INTERNAL_27 <= cpi_a_pc(28);
CPI_A_PC_INTERNAL_28 <= cpi_a_pc(29);
CPI_A_PC_INTERNAL_29 <= cpi_a_pc(30);
CPI_A_PC_INTERNAL_30 <= cpi_a_pc(31);
CPI_A_INST_INTERNAL <= cpi_a_inst(0);
CPI_A_INST_INTERNAL_0 <= cpi_a_inst(1);
CPI_A_INST_INTERNAL_1 <= cpi_a_inst(2);
CPI_A_INST_INTERNAL_2 <= cpi_a_inst(3);
CPI_A_INST_INTERNAL_3 <= cpi_a_inst(4);
CPI_A_INST_INTERNAL_4 <= cpi_a_inst(5);
CPI_A_INST_INTERNAL_5 <= cpi_a_inst(6);
CPI_A_INST_INTERNAL_6 <= cpi_a_inst(7);
CPI_A_INST_INTERNAL_7 <= cpi_a_inst(8);
CPI_A_INST_INTERNAL_8 <= cpi_a_inst(9);
CPI_A_INST_INTERNAL_9 <= cpi_a_inst(10);
CPI_A_INST_INTERNAL_10 <= cpi_a_inst(11);
CPI_A_INST_INTERNAL_11 <= cpi_a_inst(12);
CPI_A_INST_INTERNAL_12 <= cpi_a_inst(13);
CPI_A_INST_INTERNAL_13 <= cpi_a_inst(14);
CPI_A_INST_INTERNAL_14 <= cpi_a_inst(15);
CPI_A_INST_INTERNAL_15 <= cpi_a_inst(16);
CPI_A_INST_INTERNAL_16 <= cpi_a_inst(17);
CPI_A_INST_INTERNAL_17 <= cpi_a_inst(18);
CPI_A_INST_INTERNAL_18 <= cpi_a_inst(19);
CPI_A_INST_INTERNAL_19 <= cpi_a_inst(20);
CPI_A_INST_INTERNAL_20 <= cpi_a_inst(21);
CPI_A_INST_INTERNAL_21 <= cpi_a_inst(22);
CPI_A_INST_INTERNAL_22 <= cpi_a_inst(23);
CPI_A_INST_INTERNAL_23 <= cpi_a_inst(24);
CPI_A_INST_INTERNAL_24 <= cpi_a_inst(25);
CPI_A_INST_INTERNAL_25 <= cpi_a_inst(26);
CPI_A_INST_INTERNAL_26 <= cpi_a_inst(27);
CPI_A_INST_INTERNAL_27 <= cpi_a_inst(28);
CPI_A_INST_INTERNAL_28 <= cpi_a_inst(29);
CPI_A_INST_INTERNAL_29 <= cpi_a_inst(30);
CPI_A_INST_INTERNAL_30 <= cpi_a_inst(31);
CPI_A_CNT_INTERNAL <= cpi_a_cnt(0);
CPI_A_CNT_INTERNAL_0 <= cpi_a_cnt(1);
CPI_A_TRAP_INTERNAL <= cpi_a_trap;
CPI_A_ANNUL_INTERNAL <= cpi_a_annul;
CPI_A_PV_INTERNAL <= cpi_a_pv;
CPI_E_PC_INTERNAL <= cpi_e_pc(0);
CPI_E_PC_INTERNAL_0 <= cpi_e_pc(1);
CPI_E_PC_INTERNAL_1 <= cpi_e_pc(2);
CPI_E_PC_INTERNAL_2 <= cpi_e_pc(3);
CPI_E_PC_INTERNAL_3 <= cpi_e_pc(4);
CPI_E_PC_INTERNAL_4 <= cpi_e_pc(5);
CPI_E_PC_INTERNAL_5 <= cpi_e_pc(6);
CPI_E_PC_INTERNAL_6 <= cpi_e_pc(7);
CPI_E_PC_INTERNAL_7 <= cpi_e_pc(8);
CPI_E_PC_INTERNAL_8 <= cpi_e_pc(9);
CPI_E_PC_INTERNAL_9 <= cpi_e_pc(10);
CPI_E_PC_INTERNAL_10 <= cpi_e_pc(11);
CPI_E_PC_INTERNAL_11 <= cpi_e_pc(12);
CPI_E_PC_INTERNAL_12 <= cpi_e_pc(13);
CPI_E_PC_INTERNAL_13 <= cpi_e_pc(14);
CPI_E_PC_INTERNAL_14 <= cpi_e_pc(15);
CPI_E_PC_INTERNAL_15 <= cpi_e_pc(16);
CPI_E_PC_INTERNAL_16 <= cpi_e_pc(17);
CPI_E_PC_INTERNAL_17 <= cpi_e_pc(18);
CPI_E_PC_INTERNAL_18 <= cpi_e_pc(19);
CPI_E_PC_INTERNAL_19 <= cpi_e_pc(20);
CPI_E_PC_INTERNAL_20 <= cpi_e_pc(21);
CPI_E_PC_INTERNAL_21 <= cpi_e_pc(22);
CPI_E_PC_INTERNAL_22 <= cpi_e_pc(23);
CPI_E_PC_INTERNAL_23 <= cpi_e_pc(24);
CPI_E_PC_INTERNAL_24 <= cpi_e_pc(25);
CPI_E_PC_INTERNAL_25 <= cpi_e_pc(26);
CPI_E_PC_INTERNAL_26 <= cpi_e_pc(27);
CPI_E_PC_INTERNAL_27 <= cpi_e_pc(28);
CPI_E_PC_INTERNAL_28 <= cpi_e_pc(29);
CPI_E_PC_INTERNAL_29 <= cpi_e_pc(30);
CPI_E_PC_INTERNAL_30 <= cpi_e_pc(31);
CPI_E_INST_INTERNAL <= cpi_e_inst(0);
CPI_E_INST_INTERNAL_0 <= cpi_e_inst(1);
CPI_E_INST_INTERNAL_1 <= cpi_e_inst(2);
CPI_E_INST_INTERNAL_2 <= cpi_e_inst(3);
CPI_E_INST_INTERNAL_3 <= cpi_e_inst(4);
CPI_E_INST_INTERNAL_4 <= cpi_e_inst(5);
CPI_E_INST_INTERNAL_5 <= cpi_e_inst(6);
CPI_E_INST_INTERNAL_6 <= cpi_e_inst(7);
CPI_E_INST_INTERNAL_7 <= cpi_e_inst(8);
CPI_E_INST_INTERNAL_8 <= cpi_e_inst(9);
CPI_E_INST_INTERNAL_9 <= cpi_e_inst(10);
CPI_E_INST_INTERNAL_10 <= cpi_e_inst(11);
CPI_E_INST_INTERNAL_11 <= cpi_e_inst(12);
CPI_E_INST_INTERNAL_12 <= cpi_e_inst(13);
CPI_E_INST_INTERNAL_13 <= cpi_e_inst(14);
CPI_E_INST_INTERNAL_14 <= cpi_e_inst(15);
CPI_E_INST_INTERNAL_15 <= cpi_e_inst(16);
CPI_E_INST_INTERNAL_16 <= cpi_e_inst(17);
CPI_E_INST_INTERNAL_17 <= cpi_e_inst(18);
CPI_E_INST_INTERNAL_18 <= cpi_e_inst(19);
CPI_E_INST_INTERNAL_19 <= cpi_e_inst(20);
CPI_E_INST_INTERNAL_20 <= cpi_e_inst(21);
CPI_E_INST_INTERNAL_21 <= cpi_e_inst(22);
CPI_E_INST_INTERNAL_22 <= cpi_e_inst(23);
CPI_E_INST_INTERNAL_23 <= cpi_e_inst(24);
CPI_E_INST_INTERNAL_24 <= cpi_e_inst(25);
CPI_E_INST_INTERNAL_25 <= cpi_e_inst(26);
CPI_E_INST_INTERNAL_26 <= cpi_e_inst(27);
CPI_E_INST_INTERNAL_27 <= cpi_e_inst(28);
CPI_E_INST_INTERNAL_28 <= cpi_e_inst(29);
CPI_E_INST_INTERNAL_29 <= cpi_e_inst(30);
CPI_E_INST_INTERNAL_30 <= cpi_e_inst(31);
CPI_E_CNT_INTERNAL <= cpi_e_cnt(0);
CPI_E_CNT_INTERNAL_0 <= cpi_e_cnt(1);
CPI_E_TRAP_INTERNAL <= cpi_e_trap;
CPI_E_ANNUL_INTERNAL <= cpi_e_annul;
CPI_E_PV_INTERNAL <= cpi_e_pv;
CPI_M_PC_INTERNAL <= cpi_m_pc(0);
CPI_M_PC_INTERNAL_0 <= cpi_m_pc(1);
CPI_M_PC_INTERNAL_1 <= cpi_m_pc(2);
CPI_M_PC_INTERNAL_2 <= cpi_m_pc(3);
CPI_M_PC_INTERNAL_3 <= cpi_m_pc(4);
CPI_M_PC_INTERNAL_4 <= cpi_m_pc(5);
CPI_M_PC_INTERNAL_5 <= cpi_m_pc(6);
CPI_M_PC_INTERNAL_6 <= cpi_m_pc(7);
CPI_M_PC_INTERNAL_7 <= cpi_m_pc(8);
CPI_M_PC_INTERNAL_8 <= cpi_m_pc(9);
CPI_M_PC_INTERNAL_9 <= cpi_m_pc(10);
CPI_M_PC_INTERNAL_10 <= cpi_m_pc(11);
CPI_M_PC_INTERNAL_11 <= cpi_m_pc(12);
CPI_M_PC_INTERNAL_12 <= cpi_m_pc(13);
CPI_M_PC_INTERNAL_13 <= cpi_m_pc(14);
CPI_M_PC_INTERNAL_14 <= cpi_m_pc(15);
CPI_M_PC_INTERNAL_15 <= cpi_m_pc(16);
CPI_M_PC_INTERNAL_16 <= cpi_m_pc(17);
CPI_M_PC_INTERNAL_17 <= cpi_m_pc(18);
CPI_M_PC_INTERNAL_18 <= cpi_m_pc(19);
CPI_M_PC_INTERNAL_19 <= cpi_m_pc(20);
CPI_M_PC_INTERNAL_20 <= cpi_m_pc(21);
CPI_M_PC_INTERNAL_21 <= cpi_m_pc(22);
CPI_M_PC_INTERNAL_22 <= cpi_m_pc(23);
CPI_M_PC_INTERNAL_23 <= cpi_m_pc(24);
CPI_M_PC_INTERNAL_24 <= cpi_m_pc(25);
CPI_M_PC_INTERNAL_25 <= cpi_m_pc(26);
CPI_M_PC_INTERNAL_26 <= cpi_m_pc(27);
CPI_M_PC_INTERNAL_27 <= cpi_m_pc(28);
CPI_M_PC_INTERNAL_28 <= cpi_m_pc(29);
CPI_M_PC_INTERNAL_29 <= cpi_m_pc(30);
CPI_M_PC_INTERNAL_30 <= cpi_m_pc(31);
CPI_M_INST_INTERNAL <= cpi_m_inst(0);
CPI_M_INST_INTERNAL_0 <= cpi_m_inst(1);
CPI_M_INST_INTERNAL_1 <= cpi_m_inst(2);
CPI_M_INST_INTERNAL_2 <= cpi_m_inst(3);
CPI_M_INST_INTERNAL_3 <= cpi_m_inst(4);
CPI_M_INST_INTERNAL_4 <= cpi_m_inst(5);
CPI_M_INST_INTERNAL_5 <= cpi_m_inst(6);
CPI_M_INST_INTERNAL_6 <= cpi_m_inst(7);
CPI_M_INST_INTERNAL_7 <= cpi_m_inst(8);
CPI_M_INST_INTERNAL_8 <= cpi_m_inst(9);
CPI_M_INST_INTERNAL_9 <= cpi_m_inst(10);
CPI_M_INST_INTERNAL_10 <= cpi_m_inst(11);
CPI_M_INST_INTERNAL_11 <= cpi_m_inst(12);
CPI_M_INST_INTERNAL_12 <= cpi_m_inst(13);
CPI_M_INST_INTERNAL_13 <= cpi_m_inst(14);
CPI_M_INST_INTERNAL_14 <= cpi_m_inst(15);
CPI_M_INST_INTERNAL_15 <= cpi_m_inst(16);
CPI_M_INST_INTERNAL_16 <= cpi_m_inst(17);
CPI_M_INST_INTERNAL_17 <= cpi_m_inst(18);
CPI_M_INST_INTERNAL_18 <= cpi_m_inst(19);
CPI_M_INST_INTERNAL_19 <= cpi_m_inst(20);
CPI_M_INST_INTERNAL_20 <= cpi_m_inst(21);
CPI_M_INST_INTERNAL_21 <= cpi_m_inst(22);
CPI_M_INST_INTERNAL_22 <= cpi_m_inst(23);
CPI_M_INST_INTERNAL_23 <= cpi_m_inst(24);
CPI_M_INST_INTERNAL_24 <= cpi_m_inst(25);
CPI_M_INST_INTERNAL_25 <= cpi_m_inst(26);
CPI_M_INST_INTERNAL_26 <= cpi_m_inst(27);
CPI_M_INST_INTERNAL_27 <= cpi_m_inst(28);
CPI_M_INST_INTERNAL_28 <= cpi_m_inst(29);
CPI_M_INST_INTERNAL_29 <= cpi_m_inst(30);
CPI_M_INST_INTERNAL_30 <= cpi_m_inst(31);
CPI_M_CNT_INTERNAL <= cpi_m_cnt(0);
CPI_M_CNT_INTERNAL_0 <= cpi_m_cnt(1);
CPI_M_TRAP_INTERNAL <= cpi_m_trap;
CPI_M_ANNUL_INTERNAL <= cpi_m_annul;
CPI_M_PV_INTERNAL <= cpi_m_pv;
CPI_X_PC_INTERNAL <= cpi_x_pc(0);
CPI_X_PC_INTERNAL_0 <= cpi_x_pc(1);
CPI_X_PC_INTERNAL_1 <= cpi_x_pc(2);
CPI_X_PC_INTERNAL_2 <= cpi_x_pc(3);
CPI_X_PC_INTERNAL_3 <= cpi_x_pc(4);
CPI_X_PC_INTERNAL_4 <= cpi_x_pc(5);
CPI_X_PC_INTERNAL_5 <= cpi_x_pc(6);
CPI_X_PC_INTERNAL_6 <= cpi_x_pc(7);
CPI_X_PC_INTERNAL_7 <= cpi_x_pc(8);
CPI_X_PC_INTERNAL_8 <= cpi_x_pc(9);
CPI_X_PC_INTERNAL_9 <= cpi_x_pc(10);
CPI_X_PC_INTERNAL_10 <= cpi_x_pc(11);
CPI_X_PC_INTERNAL_11 <= cpi_x_pc(12);
CPI_X_PC_INTERNAL_12 <= cpi_x_pc(13);
CPI_X_PC_INTERNAL_13 <= cpi_x_pc(14);
CPI_X_PC_INTERNAL_14 <= cpi_x_pc(15);
CPI_X_PC_INTERNAL_15 <= cpi_x_pc(16);
CPI_X_PC_INTERNAL_16 <= cpi_x_pc(17);
CPI_X_PC_INTERNAL_17 <= cpi_x_pc(18);
CPI_X_PC_INTERNAL_18 <= cpi_x_pc(19);
CPI_X_PC_INTERNAL_19 <= cpi_x_pc(20);
CPI_X_PC_INTERNAL_20 <= cpi_x_pc(21);
CPI_X_PC_INTERNAL_21 <= cpi_x_pc(22);
CPI_X_PC_INTERNAL_22 <= cpi_x_pc(23);
CPI_X_PC_INTERNAL_23 <= cpi_x_pc(24);
CPI_X_PC_INTERNAL_24 <= cpi_x_pc(25);
CPI_X_PC_INTERNAL_25 <= cpi_x_pc(26);
CPI_X_PC_INTERNAL_26 <= cpi_x_pc(27);
CPI_X_PC_INTERNAL_27 <= cpi_x_pc(28);
CPI_X_PC_INTERNAL_28 <= cpi_x_pc(29);
CPI_X_PC_INTERNAL_29 <= cpi_x_pc(30);
CPI_X_PC_INTERNAL_30 <= cpi_x_pc(31);
CPI_X_INST_INTERNAL <= cpi_x_inst(0);
CPI_X_INST_INTERNAL_0 <= cpi_x_inst(1);
CPI_X_INST_INTERNAL_1 <= cpi_x_inst(2);
CPI_X_INST_INTERNAL_2 <= cpi_x_inst(3);
CPI_X_INST_INTERNAL_3 <= cpi_x_inst(4);
CPI_X_INST_INTERNAL_4 <= cpi_x_inst(5);
CPI_X_INST_INTERNAL_5 <= cpi_x_inst(6);
CPI_X_INST_INTERNAL_6 <= cpi_x_inst(7);
CPI_X_INST_INTERNAL_7 <= cpi_x_inst(8);
CPI_X_INST_INTERNAL_8 <= cpi_x_inst(9);
CPI_X_INST_INTERNAL_9 <= cpi_x_inst(10);
CPI_X_INST_INTERNAL_10 <= cpi_x_inst(11);
CPI_X_INST_INTERNAL_11 <= cpi_x_inst(12);
CPI_X_INST_INTERNAL_12 <= cpi_x_inst(13);
CPI_X_INST_INTERNAL_13 <= cpi_x_inst(14);
CPI_X_INST_INTERNAL_14 <= cpi_x_inst(15);
CPI_X_INST_INTERNAL_15 <= cpi_x_inst(16);
CPI_X_INST_INTERNAL_16 <= cpi_x_inst(17);
CPI_X_INST_INTERNAL_17 <= cpi_x_inst(18);
CPI_X_INST_INTERNAL_18 <= cpi_x_inst(19);
CPI_X_INST_INTERNAL_19 <= cpi_x_inst(20);
CPI_X_INST_INTERNAL_20 <= cpi_x_inst(21);
CPI_X_INST_INTERNAL_21 <= cpi_x_inst(22);
CPI_X_INST_INTERNAL_22 <= cpi_x_inst(23);
CPI_X_INST_INTERNAL_23 <= cpi_x_inst(24);
CPI_X_INST_INTERNAL_24 <= cpi_x_inst(25);
CPI_X_INST_INTERNAL_25 <= cpi_x_inst(26);
CPI_X_INST_INTERNAL_26 <= cpi_x_inst(27);
CPI_X_INST_INTERNAL_27 <= cpi_x_inst(28);
CPI_X_INST_INTERNAL_28 <= cpi_x_inst(29);
CPI_X_INST_INTERNAL_29 <= cpi_x_inst(30);
CPI_X_INST_INTERNAL_30 <= cpi_x_inst(31);
CPI_X_CNT_INTERNAL <= cpi_x_cnt(0);
CPI_X_CNT_INTERNAL_0 <= cpi_x_cnt(1);
CPI_X_TRAP_INTERNAL <= cpi_x_trap;
CPI_X_ANNUL_INTERNAL <= cpi_x_annul;
CPI_X_PV_INTERNAL <= cpi_x_pv;
CPI_LDDATA_INTERNAL <= cpi_lddata(0);
CPI_LDDATA_INTERNAL_0 <= cpi_lddata(1);
CPI_LDDATA_INTERNAL_1 <= cpi_lddata(2);
CPI_LDDATA_INTERNAL_2 <= cpi_lddata(3);
CPI_LDDATA_INTERNAL_3 <= cpi_lddata(4);
CPI_LDDATA_INTERNAL_4 <= cpi_lddata(5);
CPI_LDDATA_INTERNAL_5 <= cpi_lddata(6);
CPI_LDDATA_INTERNAL_6 <= cpi_lddata(7);
CPI_LDDATA_INTERNAL_7 <= cpi_lddata(8);
CPI_LDDATA_INTERNAL_8 <= cpi_lddata(9);
CPI_LDDATA_INTERNAL_9 <= cpi_lddata(10);
CPI_LDDATA_INTERNAL_10 <= cpi_lddata(11);
CPI_LDDATA_INTERNAL_11 <= cpi_lddata(12);
CPI_LDDATA_INTERNAL_12 <= cpi_lddata(13);
CPI_LDDATA_INTERNAL_13 <= cpi_lddata(14);
CPI_LDDATA_INTERNAL_14 <= cpi_lddata(15);
CPI_LDDATA_INTERNAL_15 <= cpi_lddata(16);
CPI_LDDATA_INTERNAL_16 <= cpi_lddata(17);
CPI_LDDATA_INTERNAL_17 <= cpi_lddata(18);
CPI_LDDATA_INTERNAL_18 <= cpi_lddata(19);
CPI_LDDATA_INTERNAL_19 <= cpi_lddata(20);
CPI_LDDATA_INTERNAL_20 <= cpi_lddata(21);
CPI_LDDATA_INTERNAL_21 <= cpi_lddata(22);
CPI_LDDATA_INTERNAL_22 <= cpi_lddata(23);
CPI_LDDATA_INTERNAL_23 <= cpi_lddata(24);
CPI_LDDATA_INTERNAL_24 <= cpi_lddata(25);
CPI_LDDATA_INTERNAL_25 <= cpi_lddata(26);
CPI_LDDATA_INTERNAL_26 <= cpi_lddata(27);
CPI_LDDATA_INTERNAL_27 <= cpi_lddata(28);
CPI_LDDATA_INTERNAL_28 <= cpi_lddata(29);
CPI_LDDATA_INTERNAL_29 <= cpi_lddata(30);
CPI_LDDATA_INTERNAL_30 <= cpi_lddata(31);
CPI_DBG_ENABLE_INTERNAL <= cpi_dbg_enable;
CPI_DBG_WRITE_INTERNAL <= cpi_dbg_write;
CPI_DBG_FSR_INTERNAL <= cpi_dbg_fsr;
CPI_DBG_ADDR_INTERNAL <= cpi_dbg_addr(0);
CPI_DBG_ADDR_INTERNAL_0 <= cpi_dbg_addr(1);
CPI_DBG_ADDR_INTERNAL_1 <= cpi_dbg_addr(2);
CPI_DBG_ADDR_INTERNAL_2 <= cpi_dbg_addr(3);
CPI_DBG_ADDR_INTERNAL_3 <= cpi_dbg_addr(4);
CPI_DBG_DATA_INTERNAL <= cpi_dbg_data(0);
CPI_DBG_DATA_INTERNAL_0 <= cpi_dbg_data(1);
CPI_DBG_DATA_INTERNAL_1 <= cpi_dbg_data(2);
CPI_DBG_DATA_INTERNAL_2 <= cpi_dbg_data(3);
CPI_DBG_DATA_INTERNAL_3 <= cpi_dbg_data(4);
CPI_DBG_DATA_INTERNAL_4 <= cpi_dbg_data(5);
CPI_DBG_DATA_INTERNAL_5 <= cpi_dbg_data(6);
CPI_DBG_DATA_INTERNAL_6 <= cpi_dbg_data(7);
CPI_DBG_DATA_INTERNAL_7 <= cpi_dbg_data(8);
CPI_DBG_DATA_INTERNAL_8 <= cpi_dbg_data(9);
CPI_DBG_DATA_INTERNAL_9 <= cpi_dbg_data(10);
CPI_DBG_DATA_INTERNAL_10 <= cpi_dbg_data(11);
CPI_DBG_DATA_INTERNAL_11 <= cpi_dbg_data(12);
CPI_DBG_DATA_INTERNAL_12 <= cpi_dbg_data(13);
CPI_DBG_DATA_INTERNAL_13 <= cpi_dbg_data(14);
CPI_DBG_DATA_INTERNAL_14 <= cpi_dbg_data(15);
CPI_DBG_DATA_INTERNAL_15 <= cpi_dbg_data(16);
CPI_DBG_DATA_INTERNAL_16 <= cpi_dbg_data(17);
CPI_DBG_DATA_INTERNAL_17 <= cpi_dbg_data(18);
CPI_DBG_DATA_INTERNAL_18 <= cpi_dbg_data(19);
CPI_DBG_DATA_INTERNAL_19 <= cpi_dbg_data(20);
CPI_DBG_DATA_INTERNAL_20 <= cpi_dbg_data(21);
CPI_DBG_DATA_INTERNAL_21 <= cpi_dbg_data(22);
CPI_DBG_DATA_INTERNAL_22 <= cpi_dbg_data(23);
CPI_DBG_DATA_INTERNAL_23 <= cpi_dbg_data(24);
CPI_DBG_DATA_INTERNAL_24 <= cpi_dbg_data(25);
CPI_DBG_DATA_INTERNAL_25 <= cpi_dbg_data(26);
CPI_DBG_DATA_INTERNAL_26 <= cpi_dbg_data(27);
CPI_DBG_DATA_INTERNAL_27 <= cpi_dbg_data(28);
CPI_DBG_DATA_INTERNAL_28 <= cpi_dbg_data(29);
CPI_DBG_DATA_INTERNAL_29 <= cpi_dbg_data(30);
CPI_DBG_DATA_INTERNAL_30 <= cpi_dbg_data(31);
RFO1_DATA1_INTERNAL <= rfo1_data1(0);
RFO1_DATA1_INTERNAL_0 <= rfo1_data1(1);
RFO1_DATA1_INTERNAL_1 <= rfo1_data1(2);
RFO1_DATA1_INTERNAL_2 <= rfo1_data1(3);
RFO1_DATA1_INTERNAL_3 <= rfo1_data1(4);
RFO1_DATA1_INTERNAL_4 <= rfo1_data1(5);
RFO1_DATA1_INTERNAL_5 <= rfo1_data1(6);
RFO1_DATA1_INTERNAL_6 <= rfo1_data1(7);
RFO1_DATA1_INTERNAL_7 <= rfo1_data1(8);
RFO1_DATA1_INTERNAL_8 <= rfo1_data1(9);
RFO1_DATA1_INTERNAL_9 <= rfo1_data1(10);
RFO1_DATA1_INTERNAL_10 <= rfo1_data1(11);
RFO1_DATA1_INTERNAL_11 <= rfo1_data1(12);
RFO1_DATA1_INTERNAL_12 <= rfo1_data1(13);
RFO1_DATA1_INTERNAL_13 <= rfo1_data1(14);
RFO1_DATA1_INTERNAL_14 <= rfo1_data1(15);
RFO1_DATA1_INTERNAL_15 <= rfo1_data1(16);
RFO1_DATA1_INTERNAL_16 <= rfo1_data1(17);
RFO1_DATA1_INTERNAL_17 <= rfo1_data1(18);
RFO1_DATA1_INTERNAL_18 <= rfo1_data1(19);
RFO1_DATA1_INTERNAL_19 <= rfo1_data1(20);
RFO1_DATA1_INTERNAL_20 <= rfo1_data1(21);
RFO1_DATA1_INTERNAL_21 <= rfo1_data1(22);
RFO1_DATA1_INTERNAL_22 <= rfo1_data1(23);
RFO1_DATA1_INTERNAL_23 <= rfo1_data1(24);
RFO1_DATA1_INTERNAL_24 <= rfo1_data1(25);
RFO1_DATA1_INTERNAL_25 <= rfo1_data1(26);
RFO1_DATA1_INTERNAL_26 <= rfo1_data1(27);
RFO1_DATA1_INTERNAL_27 <= rfo1_data1(28);
RFO1_DATA1_INTERNAL_28 <= rfo1_data1(29);
RFO1_DATA1_INTERNAL_29 <= rfo1_data1(30);
RFO1_DATA1_INTERNAL_30 <= rfo1_data1(31);
RFO1_DATA2_INTERNAL <= rfo1_data2(0);
RFO1_DATA2_INTERNAL_0 <= rfo1_data2(1);
RFO1_DATA2_INTERNAL_1 <= rfo1_data2(2);
RFO1_DATA2_INTERNAL_2 <= rfo1_data2(3);
RFO1_DATA2_INTERNAL_3 <= rfo1_data2(4);
RFO1_DATA2_INTERNAL_4 <= rfo1_data2(5);
RFO1_DATA2_INTERNAL_5 <= rfo1_data2(6);
RFO1_DATA2_INTERNAL_6 <= rfo1_data2(7);
RFO1_DATA2_INTERNAL_7 <= rfo1_data2(8);
RFO1_DATA2_INTERNAL_8 <= rfo1_data2(9);
RFO1_DATA2_INTERNAL_9 <= rfo1_data2(10);
RFO1_DATA2_INTERNAL_10 <= rfo1_data2(11);
RFO1_DATA2_INTERNAL_11 <= rfo1_data2(12);
RFO1_DATA2_INTERNAL_12 <= rfo1_data2(13);
RFO1_DATA2_INTERNAL_13 <= rfo1_data2(14);
RFO1_DATA2_INTERNAL_14 <= rfo1_data2(15);
RFO1_DATA2_INTERNAL_15 <= rfo1_data2(16);
RFO1_DATA2_INTERNAL_16 <= rfo1_data2(17);
RFO1_DATA2_INTERNAL_17 <= rfo1_data2(18);
RFO1_DATA2_INTERNAL_18 <= rfo1_data2(19);
RFO1_DATA2_INTERNAL_19 <= rfo1_data2(20);
RFO1_DATA2_INTERNAL_20 <= rfo1_data2(21);
RFO1_DATA2_INTERNAL_21 <= rfo1_data2(22);
RFO1_DATA2_INTERNAL_22 <= rfo1_data2(23);
RFO1_DATA2_INTERNAL_23 <= rfo1_data2(24);
RFO1_DATA2_INTERNAL_24 <= rfo1_data2(25);
RFO1_DATA2_INTERNAL_25 <= rfo1_data2(26);
RFO1_DATA2_INTERNAL_26 <= rfo1_data2(27);
RFO1_DATA2_INTERNAL_27 <= rfo1_data2(28);
RFO1_DATA2_INTERNAL_28 <= rfo1_data2(29);
RFO1_DATA2_INTERNAL_29 <= rfo1_data2(30);
RFO1_DATA2_INTERNAL_30 <= rfo1_data2(31);
RFO2_DATA1_INTERNAL <= rfo2_data1(0);
RFO2_DATA1_INTERNAL_0 <= rfo2_data1(1);
RFO2_DATA1_INTERNAL_1 <= rfo2_data1(2);
RFO2_DATA1_INTERNAL_2 <= rfo2_data1(3);
RFO2_DATA1_INTERNAL_3 <= rfo2_data1(4);
RFO2_DATA1_INTERNAL_4 <= rfo2_data1(5);
RFO2_DATA1_INTERNAL_5 <= rfo2_data1(6);
RFO2_DATA1_INTERNAL_6 <= rfo2_data1(7);
RFO2_DATA1_INTERNAL_7 <= rfo2_data1(8);
RFO2_DATA1_INTERNAL_8 <= rfo2_data1(9);
RFO2_DATA1_INTERNAL_9 <= rfo2_data1(10);
RFO2_DATA1_INTERNAL_10 <= rfo2_data1(11);
RFO2_DATA1_INTERNAL_11 <= rfo2_data1(12);
RFO2_DATA1_INTERNAL_12 <= rfo2_data1(13);
RFO2_DATA1_INTERNAL_13 <= rfo2_data1(14);
RFO2_DATA1_INTERNAL_14 <= rfo2_data1(15);
RFO2_DATA1_INTERNAL_15 <= rfo2_data1(16);
RFO2_DATA1_INTERNAL_16 <= rfo2_data1(17);
RFO2_DATA1_INTERNAL_17 <= rfo2_data1(18);
RFO2_DATA1_INTERNAL_18 <= rfo2_data1(19);
RFO2_DATA1_INTERNAL_19 <= rfo2_data1(20);
RFO2_DATA1_INTERNAL_20 <= rfo2_data1(21);
RFO2_DATA1_INTERNAL_21 <= rfo2_data1(22);
RFO2_DATA1_INTERNAL_22 <= rfo2_data1(23);
RFO2_DATA1_INTERNAL_23 <= rfo2_data1(24);
RFO2_DATA1_INTERNAL_24 <= rfo2_data1(25);
RFO2_DATA1_INTERNAL_25 <= rfo2_data1(26);
RFO2_DATA1_INTERNAL_26 <= rfo2_data1(27);
RFO2_DATA1_INTERNAL_27 <= rfo2_data1(28);
RFO2_DATA1_INTERNAL_28 <= rfo2_data1(29);
RFO2_DATA1_INTERNAL_29 <= rfo2_data1(30);
RFO2_DATA1_INTERNAL_30 <= rfo2_data1(31);
RFO2_DATA2_INTERNAL <= rfo2_data2(0);
RFO2_DATA2_INTERNAL_0 <= rfo2_data2(1);
RFO2_DATA2_INTERNAL_1 <= rfo2_data2(2);
RFO2_DATA2_INTERNAL_2 <= rfo2_data2(3);
RFO2_DATA2_INTERNAL_3 <= rfo2_data2(4);
RFO2_DATA2_INTERNAL_4 <= rfo2_data2(5);
RFO2_DATA2_INTERNAL_5 <= rfo2_data2(6);
RFO2_DATA2_INTERNAL_6 <= rfo2_data2(7);
RFO2_DATA2_INTERNAL_7 <= rfo2_data2(8);
RFO2_DATA2_INTERNAL_8 <= rfo2_data2(9);
RFO2_DATA2_INTERNAL_9 <= rfo2_data2(10);
RFO2_DATA2_INTERNAL_10 <= rfo2_data2(11);
RFO2_DATA2_INTERNAL_11 <= rfo2_data2(12);
RFO2_DATA2_INTERNAL_12 <= rfo2_data2(13);
RFO2_DATA2_INTERNAL_13 <= rfo2_data2(14);
RFO2_DATA2_INTERNAL_14 <= rfo2_data2(15);
RFO2_DATA2_INTERNAL_15 <= rfo2_data2(16);
RFO2_DATA2_INTERNAL_16 <= rfo2_data2(17);
RFO2_DATA2_INTERNAL_17 <= rfo2_data2(18);
RFO2_DATA2_INTERNAL_18 <= rfo2_data2(19);
RFO2_DATA2_INTERNAL_19 <= rfo2_data2(20);
RFO2_DATA2_INTERNAL_20 <= rfo2_data2(21);
RFO2_DATA2_INTERNAL_21 <= rfo2_data2(22);
RFO2_DATA2_INTERNAL_22 <= rfo2_data2(23);
RFO2_DATA2_INTERNAL_23 <= rfo2_data2(24);
RFO2_DATA2_INTERNAL_24 <= rfo2_data2(25);
RFO2_DATA2_INTERNAL_25 <= rfo2_data2(26);
RFO2_DATA2_INTERNAL_26 <= rfo2_data2(27);
RFO2_DATA2_INTERNAL_27 <= rfo2_data2(28);
RFO2_DATA2_INTERNAL_28 <= rfo2_data2(29);
RFO2_DATA2_INTERNAL_29 <= rfo2_data2(30);
RFO2_DATA2_INTERNAL_30 <= rfo2_data2(31);
end beh;

